/*
Copyright � 2013 lieumychuong@gmail.com

File		: 256 bit wide Crc generator
Description	:

Remarks		:

Revision	:
	Date	Author	Description

*/
module mCrc32_256(
	input [255:0] iv_Input,
	input i_SoP,
	input i_EoP,
	input i_Dv,
	input i_Clr,
	input i_Clk,
	input [4:0] i5_SoPEmpty,
	input [4:0] i5_EoPEmpty,
	output reg o_CrcV,
	output reg [31:0] o32_Crc);

	reg [31:0] r32_Crc;
	wire [31:0] w32_Crc;
	wire [31:0] w32_CrcDiv;
	reg [31:0] r32_X_n;
	reg r_End;
	
	wire [255:0] w256_LstWrdMask;
	wire [255:0] w256_FstWrdMask;
	wire [255:0] w256_In1,w256_In2;
	
	
	assign w256_In1[255:224] = r32_Crc^(iv_Input[255:224]&w256_LstWrdMask[255:224]&w256_FstWrdMask[255:224]);
	assign w256_In1[223:000] = (iv_Input[223:0]&w256_LstWrdMask[223:0]&w256_FstWrdMask[223:000]);
	
	mCrc32_256comb uCrc32(.iv_Input(w256_In1),.o32_Crc(w32_Crc));
	mGFMultiplier	uMult(.iv_PolyA(r32_Crc),.iv_PolyB(r32_X_n),.ov_PolyProd(w32_CrcDiv));
	
	generate 
		genvar I;
		for(I=0;I<32;I=I+1)
			begin:mask
			assign w256_LstWrdMask[I*8+7-:8] = (i5_EoPEmpty>I && i_EoP)?8'h00:8'hFF;
			assign w256_FstWrdMask[(32-I)*8-1-:8] = (i5_SoPEmpty>I && i_SoP)?8'h00:8'hFF;
			end		
	endgenerate
	
	always@(posedge i_Clk)
	begin 
		if(i_Clr|r_End) 
			begin 
			r32_Crc <= 32'h0;
			r32_X_n <= 32'h1;
		end
		else begin 
			if(i_Dv)  
				r32_Crc <= w32_Crc;			
		
			if(i_Dv & i_EoP)
			case(i5_EoPEmpty)
			5'd01 : r32_X_n <= 32'ha9d3e6a6;
			5'd02 : r32_X_n <= 32'h1aca48eb;
			5'd03 : r32_X_n <= 32'h876d81f8;
			5'd04 : r32_X_n <= 32'hcbf1acda;
			5'd05 : r32_X_n <= 32'hfd7384d7;
			5'd06 : r32_X_n <= 32'ha3011ff4;
			5'd07 : r32_X_n <= 32'h3c423fe9;
			5'd08 : r32_X_n <= 32'hd02dd974;
			5'd09 : r32_X_n <= 32'hbe519df4;
			5'd10 : r32_X_n <= 32'h3c5f6f6b;
			5'd11 : r32_X_n <= 32'h052b9a04;
			5'd12 : r32_X_n <= 32'haec88a6c;
			5'd13 : r32_X_n <= 32'h55c19a4a;
			5'd14 : r32_X_n <= 32'hcd39868c;
			5'd15 : r32_X_n <= 32'h753a48f0;
			5'd16 : r32_X_n <= 32'h9259a548;
			5'd17 : r32_X_n <= 32'h9a98ce48;
			5'd18 : r32_X_n <= 32'h9a900f23;
			5'd19 : r32_X_n <= 32'h9f87c289;
			5'd20 : r32_X_n <= 32'h7276b1e4;
			5'd21 : r32_X_n <= 32'h8e27f4f1;
			5'd22 : r32_X_n <= 32'h3b715e52;
			5'd23 : r32_X_n <= 32'h26b9d4a5;
			5'd24 : r32_X_n <= 32'he4f01484;
			5'd25 : r32_X_n <= 32'h2c49df39;
			5'd26 : r32_X_n <= 32'h23b9294f;
			5'd27 : r32_X_n <= 32'hca51b96f;
			5'd28 : r32_X_n <= 32'hab103524;
			5'd29 : r32_X_n <= 32'hcfced518;
			5'd30 : r32_X_n <= 32'heb212c38;
			5'd31 : r32_X_n <= 32'h8aada71a;
			default : r32_X_n <= 32'h1;
			endcase							
		end
		r_End <= i_EoP;
		o_CrcV <= r_End;
		if(r_End) 
			o32_Crc <= w32_CrcDiv;			
	end
endmodule 
	
module mGFMultiplier #(parameter pPolyOrder=31, pGenerator=32'h04C11DB7)(
	input 	[pPolyOrder:0] iv_PolyA,
	input 	[pPolyOrder:0] iv_PolyB,
	output 	[pPolyOrder:0] ov_PolyProd);
		
	wire  [pPolyOrder:0] wv_Alpha[0:pPolyOrder*2];
	wire [pPolyOrder*2:0] wv_Product;
	wire [pPolyOrder*2:0] wv_P [0:pPolyOrder*2];	
	
	generate 
		genvar I,P;
		for(I=0;I<=(pPolyOrder*2);I=I+1)
			begin:add
				for(P=0;P<=I;P=P+1)
					begin:multiply
						assign wv_P[I][P]=((P>pPolyOrder)?1'b0:iv_PolyA[P])&(((I-P)>pPolyOrder)?1'b0:iv_PolyB[I-P]); 						
					end
				assign wv_Product[I]=^wv_P[I];
			end
	endgenerate
	
	generate 
		genvar Q;
		for(Q=0;Q<(pPolyOrder*2);Q=Q+1)
		begin:zeroouttherest 
			assign wv_P[Q][pPolyOrder*2:Q+1]=0;
		end
	endgenerate
		
	assign wv_Alpha[0]=1;
	assign wv_Alpha[1]=2;
	generate 
	genvar K;
	for(K=2;K<=(pPolyOrder*2);K=K+1)
		begin:genalphak
		assign wv_Alpha[K]=(wv_Alpha[K-1][pPolyOrder])?{wv_Alpha[K-1][pPolyOrder-1:0],1'b0}^pGenerator:{wv_Alpha[K-1][pPolyOrder-1:0],1'b0};
		end
	endgenerate
	
	wire [pPolyOrder-1:0] wv_Sum [0:pPolyOrder];	
		generate 
			genvar M,N;
			for(M=0;M<=pPolyOrder;M=M+1)
				begin:row
				for(N=0;N<pPolyOrder;N=N+1)
					begin:col
						assign wv_Sum[M][N]=wv_Product[N+pPolyOrder+1]&wv_Alpha[N+pPolyOrder+1][M];						
					end	
					assign ov_PolyProd[M]=(^wv_Sum[M])^wv_Product[M];
				end
		endgenerate
endmodule


module mCrc32_256comb(
	input [255:0] iv_Input,
	output [31:0] o32_Crc);

reg [31:0] rvCrc [0:255];

always@(*)
begin
case(iv_Input[007:000])
8'h00 : rvCrc[0] <= 32'h00000000;
8'h01 : rvCrc[0] <= 32'h04c11db7;
8'h02 : rvCrc[0] <= 32'h09823b6e;
8'h03 : rvCrc[0] <= 32'h0d4326d9;
8'h04 : rvCrc[0] <= 32'h130476dc;
8'h05 : rvCrc[0] <= 32'h17c56b6b;
8'h06 : rvCrc[0] <= 32'h1a864db2;
8'h07 : rvCrc[0] <= 32'h1e475005;
8'h08 : rvCrc[0] <= 32'h2608edb8;
8'h09 : rvCrc[0] <= 32'h22c9f00f;
8'h0a : rvCrc[0] <= 32'h2f8ad6d6;
8'h0b : rvCrc[0] <= 32'h2b4bcb61;
8'h0c : rvCrc[0] <= 32'h350c9b64;
8'h0d : rvCrc[0] <= 32'h31cd86d3;
8'h0e : rvCrc[0] <= 32'h3c8ea00a;
8'h0f : rvCrc[0] <= 32'h384fbdbd;
8'h10 : rvCrc[0] <= 32'h4c11db70;
8'h11 : rvCrc[0] <= 32'h48d0c6c7;
8'h12 : rvCrc[0] <= 32'h4593e01e;
8'h13 : rvCrc[0] <= 32'h4152fda9;
8'h14 : rvCrc[0] <= 32'h5f15adac;
8'h15 : rvCrc[0] <= 32'h5bd4b01b;
8'h16 : rvCrc[0] <= 32'h569796c2;
8'h17 : rvCrc[0] <= 32'h52568b75;
8'h18 : rvCrc[0] <= 32'h6a1936c8;
8'h19 : rvCrc[0] <= 32'h6ed82b7f;
8'h1a : rvCrc[0] <= 32'h639b0da6;
8'h1b : rvCrc[0] <= 32'h675a1011;
8'h1c : rvCrc[0] <= 32'h791d4014;
8'h1d : rvCrc[0] <= 32'h7ddc5da3;
8'h1e : rvCrc[0] <= 32'h709f7b7a;
8'h1f : rvCrc[0] <= 32'h745e66cd;
8'h20 : rvCrc[0] <= 32'h9823b6e0;
8'h21 : rvCrc[0] <= 32'h9ce2ab57;
8'h22 : rvCrc[0] <= 32'h91a18d8e;
8'h23 : rvCrc[0] <= 32'h95609039;
8'h24 : rvCrc[0] <= 32'h8b27c03c;
8'h25 : rvCrc[0] <= 32'h8fe6dd8b;
8'h26 : rvCrc[0] <= 32'h82a5fb52;
8'h27 : rvCrc[0] <= 32'h8664e6e5;
8'h28 : rvCrc[0] <= 32'hbe2b5b58;
8'h29 : rvCrc[0] <= 32'hbaea46ef;
8'h2a : rvCrc[0] <= 32'hb7a96036;
8'h2b : rvCrc[0] <= 32'hb3687d81;
8'h2c : rvCrc[0] <= 32'had2f2d84;
8'h2d : rvCrc[0] <= 32'ha9ee3033;
8'h2e : rvCrc[0] <= 32'ha4ad16ea;
8'h2f : rvCrc[0] <= 32'ha06c0b5d;
8'h30 : rvCrc[0] <= 32'hd4326d90;
8'h31 : rvCrc[0] <= 32'hd0f37027;
8'h32 : rvCrc[0] <= 32'hddb056fe;
8'h33 : rvCrc[0] <= 32'hd9714b49;
8'h34 : rvCrc[0] <= 32'hc7361b4c;
8'h35 : rvCrc[0] <= 32'hc3f706fb;
8'h36 : rvCrc[0] <= 32'hceb42022;
8'h37 : rvCrc[0] <= 32'hca753d95;
8'h38 : rvCrc[0] <= 32'hf23a8028;
8'h39 : rvCrc[0] <= 32'hf6fb9d9f;
8'h3a : rvCrc[0] <= 32'hfbb8bb46;
8'h3b : rvCrc[0] <= 32'hff79a6f1;
8'h3c : rvCrc[0] <= 32'he13ef6f4;
8'h3d : rvCrc[0] <= 32'he5ffeb43;
8'h3e : rvCrc[0] <= 32'he8bccd9a;
8'h3f : rvCrc[0] <= 32'hec7dd02d;
8'h40 : rvCrc[0] <= 32'h34867077;
8'h41 : rvCrc[0] <= 32'h30476dc0;
8'h42 : rvCrc[0] <= 32'h3d044b19;
8'h43 : rvCrc[0] <= 32'h39c556ae;
8'h44 : rvCrc[0] <= 32'h278206ab;
8'h45 : rvCrc[0] <= 32'h23431b1c;
8'h46 : rvCrc[0] <= 32'h2e003dc5;
8'h47 : rvCrc[0] <= 32'h2ac12072;
8'h48 : rvCrc[0] <= 32'h128e9dcf;
8'h49 : rvCrc[0] <= 32'h164f8078;
8'h4a : rvCrc[0] <= 32'h1b0ca6a1;
8'h4b : rvCrc[0] <= 32'h1fcdbb16;
8'h4c : rvCrc[0] <= 32'h018aeb13;
8'h4d : rvCrc[0] <= 32'h054bf6a4;
8'h4e : rvCrc[0] <= 32'h0808d07d;
8'h4f : rvCrc[0] <= 32'h0cc9cdca;
8'h50 : rvCrc[0] <= 32'h7897ab07;
8'h51 : rvCrc[0] <= 32'h7c56b6b0;
8'h52 : rvCrc[0] <= 32'h71159069;
8'h53 : rvCrc[0] <= 32'h75d48dde;
8'h54 : rvCrc[0] <= 32'h6b93dddb;
8'h55 : rvCrc[0] <= 32'h6f52c06c;
8'h56 : rvCrc[0] <= 32'h6211e6b5;
8'h57 : rvCrc[0] <= 32'h66d0fb02;
8'h58 : rvCrc[0] <= 32'h5e9f46bf;
8'h59 : rvCrc[0] <= 32'h5a5e5b08;
8'h5a : rvCrc[0] <= 32'h571d7dd1;
8'h5b : rvCrc[0] <= 32'h53dc6066;
8'h5c : rvCrc[0] <= 32'h4d9b3063;
8'h5d : rvCrc[0] <= 32'h495a2dd4;
8'h5e : rvCrc[0] <= 32'h44190b0d;
8'h5f : rvCrc[0] <= 32'h40d816ba;
8'h60 : rvCrc[0] <= 32'haca5c697;
8'h61 : rvCrc[0] <= 32'ha864db20;
8'h62 : rvCrc[0] <= 32'ha527fdf9;
8'h63 : rvCrc[0] <= 32'ha1e6e04e;
8'h64 : rvCrc[0] <= 32'hbfa1b04b;
8'h65 : rvCrc[0] <= 32'hbb60adfc;
8'h66 : rvCrc[0] <= 32'hb6238b25;
8'h67 : rvCrc[0] <= 32'hb2e29692;
8'h68 : rvCrc[0] <= 32'h8aad2b2f;
8'h69 : rvCrc[0] <= 32'h8e6c3698;
8'h6a : rvCrc[0] <= 32'h832f1041;
8'h6b : rvCrc[0] <= 32'h87ee0df6;
8'h6c : rvCrc[0] <= 32'h99a95df3;
8'h6d : rvCrc[0] <= 32'h9d684044;
8'h6e : rvCrc[0] <= 32'h902b669d;
8'h6f : rvCrc[0] <= 32'h94ea7b2a;
8'h70 : rvCrc[0] <= 32'he0b41de7;
8'h71 : rvCrc[0] <= 32'he4750050;
8'h72 : rvCrc[0] <= 32'he9362689;
8'h73 : rvCrc[0] <= 32'hedf73b3e;
8'h74 : rvCrc[0] <= 32'hf3b06b3b;
8'h75 : rvCrc[0] <= 32'hf771768c;
8'h76 : rvCrc[0] <= 32'hfa325055;
8'h77 : rvCrc[0] <= 32'hfef34de2;
8'h78 : rvCrc[0] <= 32'hc6bcf05f;
8'h79 : rvCrc[0] <= 32'hc27dede8;
8'h7a : rvCrc[0] <= 32'hcf3ecb31;
8'h7b : rvCrc[0] <= 32'hcbffd686;
8'h7c : rvCrc[0] <= 32'hd5b88683;
8'h7d : rvCrc[0] <= 32'hd1799b34;
8'h7e : rvCrc[0] <= 32'hdc3abded;
8'h7f : rvCrc[0] <= 32'hd8fba05a;
8'h80 : rvCrc[0] <= 32'h690ce0ee;
8'h81 : rvCrc[0] <= 32'h6dcdfd59;
8'h82 : rvCrc[0] <= 32'h608edb80;
8'h83 : rvCrc[0] <= 32'h644fc637;
8'h84 : rvCrc[0] <= 32'h7a089632;
8'h85 : rvCrc[0] <= 32'h7ec98b85;
8'h86 : rvCrc[0] <= 32'h738aad5c;
8'h87 : rvCrc[0] <= 32'h774bb0eb;
8'h88 : rvCrc[0] <= 32'h4f040d56;
8'h89 : rvCrc[0] <= 32'h4bc510e1;
8'h8a : rvCrc[0] <= 32'h46863638;
8'h8b : rvCrc[0] <= 32'h42472b8f;
8'h8c : rvCrc[0] <= 32'h5c007b8a;
8'h8d : rvCrc[0] <= 32'h58c1663d;
8'h8e : rvCrc[0] <= 32'h558240e4;
8'h8f : rvCrc[0] <= 32'h51435d53;
8'h90 : rvCrc[0] <= 32'h251d3b9e;
8'h91 : rvCrc[0] <= 32'h21dc2629;
8'h92 : rvCrc[0] <= 32'h2c9f00f0;
8'h93 : rvCrc[0] <= 32'h285e1d47;
8'h94 : rvCrc[0] <= 32'h36194d42;
8'h95 : rvCrc[0] <= 32'h32d850f5;
8'h96 : rvCrc[0] <= 32'h3f9b762c;
8'h97 : rvCrc[0] <= 32'h3b5a6b9b;
8'h98 : rvCrc[0] <= 32'h0315d626;
8'h99 : rvCrc[0] <= 32'h07d4cb91;
8'h9a : rvCrc[0] <= 32'h0a97ed48;
8'h9b : rvCrc[0] <= 32'h0e56f0ff;
8'h9c : rvCrc[0] <= 32'h1011a0fa;
8'h9d : rvCrc[0] <= 32'h14d0bd4d;
8'h9e : rvCrc[0] <= 32'h19939b94;
8'h9f : rvCrc[0] <= 32'h1d528623;
8'ha0 : rvCrc[0] <= 32'hf12f560e;
8'ha1 : rvCrc[0] <= 32'hf5ee4bb9;
8'ha2 : rvCrc[0] <= 32'hf8ad6d60;
8'ha3 : rvCrc[0] <= 32'hfc6c70d7;
8'ha4 : rvCrc[0] <= 32'he22b20d2;
8'ha5 : rvCrc[0] <= 32'he6ea3d65;
8'ha6 : rvCrc[0] <= 32'heba91bbc;
8'ha7 : rvCrc[0] <= 32'hef68060b;
8'ha8 : rvCrc[0] <= 32'hd727bbb6;
8'ha9 : rvCrc[0] <= 32'hd3e6a601;
8'haa : rvCrc[0] <= 32'hdea580d8;
8'hab : rvCrc[0] <= 32'hda649d6f;
8'hac : rvCrc[0] <= 32'hc423cd6a;
8'had : rvCrc[0] <= 32'hc0e2d0dd;
8'hae : rvCrc[0] <= 32'hcda1f604;
8'haf : rvCrc[0] <= 32'hc960ebb3;
8'hb0 : rvCrc[0] <= 32'hbd3e8d7e;
8'hb1 : rvCrc[0] <= 32'hb9ff90c9;
8'hb2 : rvCrc[0] <= 32'hb4bcb610;
8'hb3 : rvCrc[0] <= 32'hb07daba7;
8'hb4 : rvCrc[0] <= 32'hae3afba2;
8'hb5 : rvCrc[0] <= 32'haafbe615;
8'hb6 : rvCrc[0] <= 32'ha7b8c0cc;
8'hb7 : rvCrc[0] <= 32'ha379dd7b;
8'hb8 : rvCrc[0] <= 32'h9b3660c6;
8'hb9 : rvCrc[0] <= 32'h9ff77d71;
8'hba : rvCrc[0] <= 32'h92b45ba8;
8'hbb : rvCrc[0] <= 32'h9675461f;
8'hbc : rvCrc[0] <= 32'h8832161a;
8'hbd : rvCrc[0] <= 32'h8cf30bad;
8'hbe : rvCrc[0] <= 32'h81b02d74;
8'hbf : rvCrc[0] <= 32'h857130c3;
8'hc0 : rvCrc[0] <= 32'h5d8a9099;
8'hc1 : rvCrc[0] <= 32'h594b8d2e;
8'hc2 : rvCrc[0] <= 32'h5408abf7;
8'hc3 : rvCrc[0] <= 32'h50c9b640;
8'hc4 : rvCrc[0] <= 32'h4e8ee645;
8'hc5 : rvCrc[0] <= 32'h4a4ffbf2;
8'hc6 : rvCrc[0] <= 32'h470cdd2b;
8'hc7 : rvCrc[0] <= 32'h43cdc09c;
8'hc8 : rvCrc[0] <= 32'h7b827d21;
8'hc9 : rvCrc[0] <= 32'h7f436096;
8'hca : rvCrc[0] <= 32'h7200464f;
8'hcb : rvCrc[0] <= 32'h76c15bf8;
8'hcc : rvCrc[0] <= 32'h68860bfd;
8'hcd : rvCrc[0] <= 32'h6c47164a;
8'hce : rvCrc[0] <= 32'h61043093;
8'hcf : rvCrc[0] <= 32'h65c52d24;
8'hd0 : rvCrc[0] <= 32'h119b4be9;
8'hd1 : rvCrc[0] <= 32'h155a565e;
8'hd2 : rvCrc[0] <= 32'h18197087;
8'hd3 : rvCrc[0] <= 32'h1cd86d30;
8'hd4 : rvCrc[0] <= 32'h029f3d35;
8'hd5 : rvCrc[0] <= 32'h065e2082;
8'hd6 : rvCrc[0] <= 32'h0b1d065b;
8'hd7 : rvCrc[0] <= 32'h0fdc1bec;
8'hd8 : rvCrc[0] <= 32'h3793a651;
8'hd9 : rvCrc[0] <= 32'h3352bbe6;
8'hda : rvCrc[0] <= 32'h3e119d3f;
8'hdb : rvCrc[0] <= 32'h3ad08088;
8'hdc : rvCrc[0] <= 32'h2497d08d;
8'hdd : rvCrc[0] <= 32'h2056cd3a;
8'hde : rvCrc[0] <= 32'h2d15ebe3;
8'hdf : rvCrc[0] <= 32'h29d4f654;
8'he0 : rvCrc[0] <= 32'hc5a92679;
8'he1 : rvCrc[0] <= 32'hc1683bce;
8'he2 : rvCrc[0] <= 32'hcc2b1d17;
8'he3 : rvCrc[0] <= 32'hc8ea00a0;
8'he4 : rvCrc[0] <= 32'hd6ad50a5;
8'he5 : rvCrc[0] <= 32'hd26c4d12;
8'he6 : rvCrc[0] <= 32'hdf2f6bcb;
8'he7 : rvCrc[0] <= 32'hdbee767c;
8'he8 : rvCrc[0] <= 32'he3a1cbc1;
8'he9 : rvCrc[0] <= 32'he760d676;
8'hea : rvCrc[0] <= 32'hea23f0af;
8'heb : rvCrc[0] <= 32'heee2ed18;
8'hec : rvCrc[0] <= 32'hf0a5bd1d;
8'hed : rvCrc[0] <= 32'hf464a0aa;
8'hee : rvCrc[0] <= 32'hf9278673;
8'hef : rvCrc[0] <= 32'hfde69bc4;
8'hf0 : rvCrc[0] <= 32'h89b8fd09;
8'hf1 : rvCrc[0] <= 32'h8d79e0be;
8'hf2 : rvCrc[0] <= 32'h803ac667;
8'hf3 : rvCrc[0] <= 32'h84fbdbd0;
8'hf4 : rvCrc[0] <= 32'h9abc8bd5;
8'hf5 : rvCrc[0] <= 32'h9e7d9662;
8'hf6 : rvCrc[0] <= 32'h933eb0bb;
8'hf7 : rvCrc[0] <= 32'h97ffad0c;
8'hf8 : rvCrc[0] <= 32'hafb010b1;
8'hf9 : rvCrc[0] <= 32'hab710d06;
8'hfa : rvCrc[0] <= 32'ha6322bdf;
8'hfb : rvCrc[0] <= 32'ha2f33668;
8'hfc : rvCrc[0] <= 32'hbcb4666d;
8'hfd : rvCrc[0] <= 32'hb8757bda;
8'hfe : rvCrc[0] <= 32'hb5365d03;
8'hff : rvCrc[0] <= 32'hb1f740b4;
endcase
case(iv_Input[015:008])
8'h00 : rvCrc[1] <= 32'h00000000;
8'h01 : rvCrc[1] <= 32'hd219c1dc;
8'h02 : rvCrc[1] <= 32'ha0f29e0f;
8'h03 : rvCrc[1] <= 32'h72eb5fd3;
8'h04 : rvCrc[1] <= 32'h452421a9;
8'h05 : rvCrc[1] <= 32'h973de075;
8'h06 : rvCrc[1] <= 32'he5d6bfa6;
8'h07 : rvCrc[1] <= 32'h37cf7e7a;
8'h08 : rvCrc[1] <= 32'h8a484352;
8'h09 : rvCrc[1] <= 32'h5851828e;
8'h0a : rvCrc[1] <= 32'h2abadd5d;
8'h0b : rvCrc[1] <= 32'hf8a31c81;
8'h0c : rvCrc[1] <= 32'hcf6c62fb;
8'h0d : rvCrc[1] <= 32'h1d75a327;
8'h0e : rvCrc[1] <= 32'h6f9efcf4;
8'h0f : rvCrc[1] <= 32'hbd873d28;
8'h10 : rvCrc[1] <= 32'h10519b13;
8'h11 : rvCrc[1] <= 32'hc2485acf;
8'h12 : rvCrc[1] <= 32'hb0a3051c;
8'h13 : rvCrc[1] <= 32'h62bac4c0;
8'h14 : rvCrc[1] <= 32'h5575baba;
8'h15 : rvCrc[1] <= 32'h876c7b66;
8'h16 : rvCrc[1] <= 32'hf58724b5;
8'h17 : rvCrc[1] <= 32'h279ee569;
8'h18 : rvCrc[1] <= 32'h9a19d841;
8'h19 : rvCrc[1] <= 32'h4800199d;
8'h1a : rvCrc[1] <= 32'h3aeb464e;
8'h1b : rvCrc[1] <= 32'he8f28792;
8'h1c : rvCrc[1] <= 32'hdf3df9e8;
8'h1d : rvCrc[1] <= 32'h0d243834;
8'h1e : rvCrc[1] <= 32'h7fcf67e7;
8'h1f : rvCrc[1] <= 32'hadd6a63b;
8'h20 : rvCrc[1] <= 32'h20a33626;
8'h21 : rvCrc[1] <= 32'hf2baf7fa;
8'h22 : rvCrc[1] <= 32'h8051a829;
8'h23 : rvCrc[1] <= 32'h524869f5;
8'h24 : rvCrc[1] <= 32'h6587178f;
8'h25 : rvCrc[1] <= 32'hb79ed653;
8'h26 : rvCrc[1] <= 32'hc5758980;
8'h27 : rvCrc[1] <= 32'h176c485c;
8'h28 : rvCrc[1] <= 32'haaeb7574;
8'h29 : rvCrc[1] <= 32'h78f2b4a8;
8'h2a : rvCrc[1] <= 32'h0a19eb7b;
8'h2b : rvCrc[1] <= 32'hd8002aa7;
8'h2c : rvCrc[1] <= 32'hefcf54dd;
8'h2d : rvCrc[1] <= 32'h3dd69501;
8'h2e : rvCrc[1] <= 32'h4f3dcad2;
8'h2f : rvCrc[1] <= 32'h9d240b0e;
8'h30 : rvCrc[1] <= 32'h30f2ad35;
8'h31 : rvCrc[1] <= 32'he2eb6ce9;
8'h32 : rvCrc[1] <= 32'h9000333a;
8'h33 : rvCrc[1] <= 32'h4219f2e6;
8'h34 : rvCrc[1] <= 32'h75d68c9c;
8'h35 : rvCrc[1] <= 32'ha7cf4d40;
8'h36 : rvCrc[1] <= 32'hd5241293;
8'h37 : rvCrc[1] <= 32'h073dd34f;
8'h38 : rvCrc[1] <= 32'hbabaee67;
8'h39 : rvCrc[1] <= 32'h68a32fbb;
8'h3a : rvCrc[1] <= 32'h1a487068;
8'h3b : rvCrc[1] <= 32'hc851b1b4;
8'h3c : rvCrc[1] <= 32'hff9ecfce;
8'h3d : rvCrc[1] <= 32'h2d870e12;
8'h3e : rvCrc[1] <= 32'h5f6c51c1;
8'h3f : rvCrc[1] <= 32'h8d75901d;
8'h40 : rvCrc[1] <= 32'h41466c4c;
8'h41 : rvCrc[1] <= 32'h935fad90;
8'h42 : rvCrc[1] <= 32'he1b4f243;
8'h43 : rvCrc[1] <= 32'h33ad339f;
8'h44 : rvCrc[1] <= 32'h04624de5;
8'h45 : rvCrc[1] <= 32'hd67b8c39;
8'h46 : rvCrc[1] <= 32'ha490d3ea;
8'h47 : rvCrc[1] <= 32'h76891236;
8'h48 : rvCrc[1] <= 32'hcb0e2f1e;
8'h49 : rvCrc[1] <= 32'h1917eec2;
8'h4a : rvCrc[1] <= 32'h6bfcb111;
8'h4b : rvCrc[1] <= 32'hb9e570cd;
8'h4c : rvCrc[1] <= 32'h8e2a0eb7;
8'h4d : rvCrc[1] <= 32'h5c33cf6b;
8'h4e : rvCrc[1] <= 32'h2ed890b8;
8'h4f : rvCrc[1] <= 32'hfcc15164;
8'h50 : rvCrc[1] <= 32'h5117f75f;
8'h51 : rvCrc[1] <= 32'h830e3683;
8'h52 : rvCrc[1] <= 32'hf1e56950;
8'h53 : rvCrc[1] <= 32'h23fca88c;
8'h54 : rvCrc[1] <= 32'h1433d6f6;
8'h55 : rvCrc[1] <= 32'hc62a172a;
8'h56 : rvCrc[1] <= 32'hb4c148f9;
8'h57 : rvCrc[1] <= 32'h66d88925;
8'h58 : rvCrc[1] <= 32'hdb5fb40d;
8'h59 : rvCrc[1] <= 32'h094675d1;
8'h5a : rvCrc[1] <= 32'h7bad2a02;
8'h5b : rvCrc[1] <= 32'ha9b4ebde;
8'h5c : rvCrc[1] <= 32'h9e7b95a4;
8'h5d : rvCrc[1] <= 32'h4c625478;
8'h5e : rvCrc[1] <= 32'h3e890bab;
8'h5f : rvCrc[1] <= 32'hec90ca77;
8'h60 : rvCrc[1] <= 32'h61e55a6a;
8'h61 : rvCrc[1] <= 32'hb3fc9bb6;
8'h62 : rvCrc[1] <= 32'hc117c465;
8'h63 : rvCrc[1] <= 32'h130e05b9;
8'h64 : rvCrc[1] <= 32'h24c17bc3;
8'h65 : rvCrc[1] <= 32'hf6d8ba1f;
8'h66 : rvCrc[1] <= 32'h8433e5cc;
8'h67 : rvCrc[1] <= 32'h562a2410;
8'h68 : rvCrc[1] <= 32'hebad1938;
8'h69 : rvCrc[1] <= 32'h39b4d8e4;
8'h6a : rvCrc[1] <= 32'h4b5f8737;
8'h6b : rvCrc[1] <= 32'h994646eb;
8'h6c : rvCrc[1] <= 32'hae893891;
8'h6d : rvCrc[1] <= 32'h7c90f94d;
8'h6e : rvCrc[1] <= 32'h0e7ba69e;
8'h6f : rvCrc[1] <= 32'hdc626742;
8'h70 : rvCrc[1] <= 32'h71b4c179;
8'h71 : rvCrc[1] <= 32'ha3ad00a5;
8'h72 : rvCrc[1] <= 32'hd1465f76;
8'h73 : rvCrc[1] <= 32'h035f9eaa;
8'h74 : rvCrc[1] <= 32'h3490e0d0;
8'h75 : rvCrc[1] <= 32'he689210c;
8'h76 : rvCrc[1] <= 32'h94627edf;
8'h77 : rvCrc[1] <= 32'h467bbf03;
8'h78 : rvCrc[1] <= 32'hfbfc822b;
8'h79 : rvCrc[1] <= 32'h29e543f7;
8'h7a : rvCrc[1] <= 32'h5b0e1c24;
8'h7b : rvCrc[1] <= 32'h8917ddf8;
8'h7c : rvCrc[1] <= 32'hbed8a382;
8'h7d : rvCrc[1] <= 32'h6cc1625e;
8'h7e : rvCrc[1] <= 32'h1e2a3d8d;
8'h7f : rvCrc[1] <= 32'hcc33fc51;
8'h80 : rvCrc[1] <= 32'h828cd898;
8'h81 : rvCrc[1] <= 32'h50951944;
8'h82 : rvCrc[1] <= 32'h227e4697;
8'h83 : rvCrc[1] <= 32'hf067874b;
8'h84 : rvCrc[1] <= 32'hc7a8f931;
8'h85 : rvCrc[1] <= 32'h15b138ed;
8'h86 : rvCrc[1] <= 32'h675a673e;
8'h87 : rvCrc[1] <= 32'hb543a6e2;
8'h88 : rvCrc[1] <= 32'h08c49bca;
8'h89 : rvCrc[1] <= 32'hdadd5a16;
8'h8a : rvCrc[1] <= 32'ha83605c5;
8'h8b : rvCrc[1] <= 32'h7a2fc419;
8'h8c : rvCrc[1] <= 32'h4de0ba63;
8'h8d : rvCrc[1] <= 32'h9ff97bbf;
8'h8e : rvCrc[1] <= 32'hed12246c;
8'h8f : rvCrc[1] <= 32'h3f0be5b0;
8'h90 : rvCrc[1] <= 32'h92dd438b;
8'h91 : rvCrc[1] <= 32'h40c48257;
8'h92 : rvCrc[1] <= 32'h322fdd84;
8'h93 : rvCrc[1] <= 32'he0361c58;
8'h94 : rvCrc[1] <= 32'hd7f96222;
8'h95 : rvCrc[1] <= 32'h05e0a3fe;
8'h96 : rvCrc[1] <= 32'h770bfc2d;
8'h97 : rvCrc[1] <= 32'ha5123df1;
8'h98 : rvCrc[1] <= 32'h189500d9;
8'h99 : rvCrc[1] <= 32'hca8cc105;
8'h9a : rvCrc[1] <= 32'hb8679ed6;
8'h9b : rvCrc[1] <= 32'h6a7e5f0a;
8'h9c : rvCrc[1] <= 32'h5db12170;
8'h9d : rvCrc[1] <= 32'h8fa8e0ac;
8'h9e : rvCrc[1] <= 32'hfd43bf7f;
8'h9f : rvCrc[1] <= 32'h2f5a7ea3;
8'ha0 : rvCrc[1] <= 32'ha22feebe;
8'ha1 : rvCrc[1] <= 32'h70362f62;
8'ha2 : rvCrc[1] <= 32'h02dd70b1;
8'ha3 : rvCrc[1] <= 32'hd0c4b16d;
8'ha4 : rvCrc[1] <= 32'he70bcf17;
8'ha5 : rvCrc[1] <= 32'h35120ecb;
8'ha6 : rvCrc[1] <= 32'h47f95118;
8'ha7 : rvCrc[1] <= 32'h95e090c4;
8'ha8 : rvCrc[1] <= 32'h2867adec;
8'ha9 : rvCrc[1] <= 32'hfa7e6c30;
8'haa : rvCrc[1] <= 32'h889533e3;
8'hab : rvCrc[1] <= 32'h5a8cf23f;
8'hac : rvCrc[1] <= 32'h6d438c45;
8'had : rvCrc[1] <= 32'hbf5a4d99;
8'hae : rvCrc[1] <= 32'hcdb1124a;
8'haf : rvCrc[1] <= 32'h1fa8d396;
8'hb0 : rvCrc[1] <= 32'hb27e75ad;
8'hb1 : rvCrc[1] <= 32'h6067b471;
8'hb2 : rvCrc[1] <= 32'h128ceba2;
8'hb3 : rvCrc[1] <= 32'hc0952a7e;
8'hb4 : rvCrc[1] <= 32'hf75a5404;
8'hb5 : rvCrc[1] <= 32'h254395d8;
8'hb6 : rvCrc[1] <= 32'h57a8ca0b;
8'hb7 : rvCrc[1] <= 32'h85b10bd7;
8'hb8 : rvCrc[1] <= 32'h383636ff;
8'hb9 : rvCrc[1] <= 32'hea2ff723;
8'hba : rvCrc[1] <= 32'h98c4a8f0;
8'hbb : rvCrc[1] <= 32'h4add692c;
8'hbc : rvCrc[1] <= 32'h7d121756;
8'hbd : rvCrc[1] <= 32'haf0bd68a;
8'hbe : rvCrc[1] <= 32'hdde08959;
8'hbf : rvCrc[1] <= 32'h0ff94885;
8'hc0 : rvCrc[1] <= 32'hc3cab4d4;
8'hc1 : rvCrc[1] <= 32'h11d37508;
8'hc2 : rvCrc[1] <= 32'h63382adb;
8'hc3 : rvCrc[1] <= 32'hb121eb07;
8'hc4 : rvCrc[1] <= 32'h86ee957d;
8'hc5 : rvCrc[1] <= 32'h54f754a1;
8'hc6 : rvCrc[1] <= 32'h261c0b72;
8'hc7 : rvCrc[1] <= 32'hf405caae;
8'hc8 : rvCrc[1] <= 32'h4982f786;
8'hc9 : rvCrc[1] <= 32'h9b9b365a;
8'hca : rvCrc[1] <= 32'he9706989;
8'hcb : rvCrc[1] <= 32'h3b69a855;
8'hcc : rvCrc[1] <= 32'h0ca6d62f;
8'hcd : rvCrc[1] <= 32'hdebf17f3;
8'hce : rvCrc[1] <= 32'hac544820;
8'hcf : rvCrc[1] <= 32'h7e4d89fc;
8'hd0 : rvCrc[1] <= 32'hd39b2fc7;
8'hd1 : rvCrc[1] <= 32'h0182ee1b;
8'hd2 : rvCrc[1] <= 32'h7369b1c8;
8'hd3 : rvCrc[1] <= 32'ha1707014;
8'hd4 : rvCrc[1] <= 32'h96bf0e6e;
8'hd5 : rvCrc[1] <= 32'h44a6cfb2;
8'hd6 : rvCrc[1] <= 32'h364d9061;
8'hd7 : rvCrc[1] <= 32'he45451bd;
8'hd8 : rvCrc[1] <= 32'h59d36c95;
8'hd9 : rvCrc[1] <= 32'h8bcaad49;
8'hda : rvCrc[1] <= 32'hf921f29a;
8'hdb : rvCrc[1] <= 32'h2b383346;
8'hdc : rvCrc[1] <= 32'h1cf74d3c;
8'hdd : rvCrc[1] <= 32'hceee8ce0;
8'hde : rvCrc[1] <= 32'hbc05d333;
8'hdf : rvCrc[1] <= 32'h6e1c12ef;
8'he0 : rvCrc[1] <= 32'he36982f2;
8'he1 : rvCrc[1] <= 32'h3170432e;
8'he2 : rvCrc[1] <= 32'h439b1cfd;
8'he3 : rvCrc[1] <= 32'h9182dd21;
8'he4 : rvCrc[1] <= 32'ha64da35b;
8'he5 : rvCrc[1] <= 32'h74546287;
8'he6 : rvCrc[1] <= 32'h06bf3d54;
8'he7 : rvCrc[1] <= 32'hd4a6fc88;
8'he8 : rvCrc[1] <= 32'h6921c1a0;
8'he9 : rvCrc[1] <= 32'hbb38007c;
8'hea : rvCrc[1] <= 32'hc9d35faf;
8'heb : rvCrc[1] <= 32'h1bca9e73;
8'hec : rvCrc[1] <= 32'h2c05e009;
8'hed : rvCrc[1] <= 32'hfe1c21d5;
8'hee : rvCrc[1] <= 32'h8cf77e06;
8'hef : rvCrc[1] <= 32'h5eeebfda;
8'hf0 : rvCrc[1] <= 32'hf33819e1;
8'hf1 : rvCrc[1] <= 32'h2121d83d;
8'hf2 : rvCrc[1] <= 32'h53ca87ee;
8'hf3 : rvCrc[1] <= 32'h81d34632;
8'hf4 : rvCrc[1] <= 32'hb61c3848;
8'hf5 : rvCrc[1] <= 32'h6405f994;
8'hf6 : rvCrc[1] <= 32'h16eea647;
8'hf7 : rvCrc[1] <= 32'hc4f7679b;
8'hf8 : rvCrc[1] <= 32'h79705ab3;
8'hf9 : rvCrc[1] <= 32'hab699b6f;
8'hfa : rvCrc[1] <= 32'hd982c4bc;
8'hfb : rvCrc[1] <= 32'h0b9b0560;
8'hfc : rvCrc[1] <= 32'h3c547b1a;
8'hfd : rvCrc[1] <= 32'hee4dbac6;
8'hfe : rvCrc[1] <= 32'h9ca6e515;
8'hff : rvCrc[1] <= 32'h4ebf24c9;
endcase
case(iv_Input[023:016])
8'h00 : rvCrc[2] <= 32'h00000000;
8'h01 : rvCrc[2] <= 32'h01d8ac87;
8'h02 : rvCrc[2] <= 32'h03b1590e;
8'h03 : rvCrc[2] <= 32'h0269f589;
8'h04 : rvCrc[2] <= 32'h0762b21c;
8'h05 : rvCrc[2] <= 32'h06ba1e9b;
8'h06 : rvCrc[2] <= 32'h04d3eb12;
8'h07 : rvCrc[2] <= 32'h050b4795;
8'h08 : rvCrc[2] <= 32'h0ec56438;
8'h09 : rvCrc[2] <= 32'h0f1dc8bf;
8'h0a : rvCrc[2] <= 32'h0d743d36;
8'h0b : rvCrc[2] <= 32'h0cac91b1;
8'h0c : rvCrc[2] <= 32'h09a7d624;
8'h0d : rvCrc[2] <= 32'h087f7aa3;
8'h0e : rvCrc[2] <= 32'h0a168f2a;
8'h0f : rvCrc[2] <= 32'h0bce23ad;
8'h10 : rvCrc[2] <= 32'h1d8ac870;
8'h11 : rvCrc[2] <= 32'h1c5264f7;
8'h12 : rvCrc[2] <= 32'h1e3b917e;
8'h13 : rvCrc[2] <= 32'h1fe33df9;
8'h14 : rvCrc[2] <= 32'h1ae87a6c;
8'h15 : rvCrc[2] <= 32'h1b30d6eb;
8'h16 : rvCrc[2] <= 32'h19592362;
8'h17 : rvCrc[2] <= 32'h18818fe5;
8'h18 : rvCrc[2] <= 32'h134fac48;
8'h19 : rvCrc[2] <= 32'h129700cf;
8'h1a : rvCrc[2] <= 32'h10fef546;
8'h1b : rvCrc[2] <= 32'h112659c1;
8'h1c : rvCrc[2] <= 32'h142d1e54;
8'h1d : rvCrc[2] <= 32'h15f5b2d3;
8'h1e : rvCrc[2] <= 32'h179c475a;
8'h1f : rvCrc[2] <= 32'h1644ebdd;
8'h20 : rvCrc[2] <= 32'h3b1590e0;
8'h21 : rvCrc[2] <= 32'h3acd3c67;
8'h22 : rvCrc[2] <= 32'h38a4c9ee;
8'h23 : rvCrc[2] <= 32'h397c6569;
8'h24 : rvCrc[2] <= 32'h3c7722fc;
8'h25 : rvCrc[2] <= 32'h3daf8e7b;
8'h26 : rvCrc[2] <= 32'h3fc67bf2;
8'h27 : rvCrc[2] <= 32'h3e1ed775;
8'h28 : rvCrc[2] <= 32'h35d0f4d8;
8'h29 : rvCrc[2] <= 32'h3408585f;
8'h2a : rvCrc[2] <= 32'h3661add6;
8'h2b : rvCrc[2] <= 32'h37b90151;
8'h2c : rvCrc[2] <= 32'h32b246c4;
8'h2d : rvCrc[2] <= 32'h336aea43;
8'h2e : rvCrc[2] <= 32'h31031fca;
8'h2f : rvCrc[2] <= 32'h30dbb34d;
8'h30 : rvCrc[2] <= 32'h269f5890;
8'h31 : rvCrc[2] <= 32'h2747f417;
8'h32 : rvCrc[2] <= 32'h252e019e;
8'h33 : rvCrc[2] <= 32'h24f6ad19;
8'h34 : rvCrc[2] <= 32'h21fdea8c;
8'h35 : rvCrc[2] <= 32'h2025460b;
8'h36 : rvCrc[2] <= 32'h224cb382;
8'h37 : rvCrc[2] <= 32'h23941f05;
8'h38 : rvCrc[2] <= 32'h285a3ca8;
8'h39 : rvCrc[2] <= 32'h2982902f;
8'h3a : rvCrc[2] <= 32'h2beb65a6;
8'h3b : rvCrc[2] <= 32'h2a33c921;
8'h3c : rvCrc[2] <= 32'h2f388eb4;
8'h3d : rvCrc[2] <= 32'h2ee02233;
8'h3e : rvCrc[2] <= 32'h2c89d7ba;
8'h3f : rvCrc[2] <= 32'h2d517b3d;
8'h40 : rvCrc[2] <= 32'h762b21c0;
8'h41 : rvCrc[2] <= 32'h77f38d47;
8'h42 : rvCrc[2] <= 32'h759a78ce;
8'h43 : rvCrc[2] <= 32'h7442d449;
8'h44 : rvCrc[2] <= 32'h714993dc;
8'h45 : rvCrc[2] <= 32'h70913f5b;
8'h46 : rvCrc[2] <= 32'h72f8cad2;
8'h47 : rvCrc[2] <= 32'h73206655;
8'h48 : rvCrc[2] <= 32'h78ee45f8;
8'h49 : rvCrc[2] <= 32'h7936e97f;
8'h4a : rvCrc[2] <= 32'h7b5f1cf6;
8'h4b : rvCrc[2] <= 32'h7a87b071;
8'h4c : rvCrc[2] <= 32'h7f8cf7e4;
8'h4d : rvCrc[2] <= 32'h7e545b63;
8'h4e : rvCrc[2] <= 32'h7c3daeea;
8'h4f : rvCrc[2] <= 32'h7de5026d;
8'h50 : rvCrc[2] <= 32'h6ba1e9b0;
8'h51 : rvCrc[2] <= 32'h6a794537;
8'h52 : rvCrc[2] <= 32'h6810b0be;
8'h53 : rvCrc[2] <= 32'h69c81c39;
8'h54 : rvCrc[2] <= 32'h6cc35bac;
8'h55 : rvCrc[2] <= 32'h6d1bf72b;
8'h56 : rvCrc[2] <= 32'h6f7202a2;
8'h57 : rvCrc[2] <= 32'h6eaaae25;
8'h58 : rvCrc[2] <= 32'h65648d88;
8'h59 : rvCrc[2] <= 32'h64bc210f;
8'h5a : rvCrc[2] <= 32'h66d5d486;
8'h5b : rvCrc[2] <= 32'h670d7801;
8'h5c : rvCrc[2] <= 32'h62063f94;
8'h5d : rvCrc[2] <= 32'h63de9313;
8'h5e : rvCrc[2] <= 32'h61b7669a;
8'h5f : rvCrc[2] <= 32'h606fca1d;
8'h60 : rvCrc[2] <= 32'h4d3eb120;
8'h61 : rvCrc[2] <= 32'h4ce61da7;
8'h62 : rvCrc[2] <= 32'h4e8fe82e;
8'h63 : rvCrc[2] <= 32'h4f5744a9;
8'h64 : rvCrc[2] <= 32'h4a5c033c;
8'h65 : rvCrc[2] <= 32'h4b84afbb;
8'h66 : rvCrc[2] <= 32'h49ed5a32;
8'h67 : rvCrc[2] <= 32'h4835f6b5;
8'h68 : rvCrc[2] <= 32'h43fbd518;
8'h69 : rvCrc[2] <= 32'h4223799f;
8'h6a : rvCrc[2] <= 32'h404a8c16;
8'h6b : rvCrc[2] <= 32'h41922091;
8'h6c : rvCrc[2] <= 32'h44996704;
8'h6d : rvCrc[2] <= 32'h4541cb83;
8'h6e : rvCrc[2] <= 32'h47283e0a;
8'h6f : rvCrc[2] <= 32'h46f0928d;
8'h70 : rvCrc[2] <= 32'h50b47950;
8'h71 : rvCrc[2] <= 32'h516cd5d7;
8'h72 : rvCrc[2] <= 32'h5305205e;
8'h73 : rvCrc[2] <= 32'h52dd8cd9;
8'h74 : rvCrc[2] <= 32'h57d6cb4c;
8'h75 : rvCrc[2] <= 32'h560e67cb;
8'h76 : rvCrc[2] <= 32'h54679242;
8'h77 : rvCrc[2] <= 32'h55bf3ec5;
8'h78 : rvCrc[2] <= 32'h5e711d68;
8'h79 : rvCrc[2] <= 32'h5fa9b1ef;
8'h7a : rvCrc[2] <= 32'h5dc04466;
8'h7b : rvCrc[2] <= 32'h5c18e8e1;
8'h7c : rvCrc[2] <= 32'h5913af74;
8'h7d : rvCrc[2] <= 32'h58cb03f3;
8'h7e : rvCrc[2] <= 32'h5aa2f67a;
8'h7f : rvCrc[2] <= 32'h5b7a5afd;
8'h80 : rvCrc[2] <= 32'hec564380;
8'h81 : rvCrc[2] <= 32'hed8eef07;
8'h82 : rvCrc[2] <= 32'hefe71a8e;
8'h83 : rvCrc[2] <= 32'hee3fb609;
8'h84 : rvCrc[2] <= 32'heb34f19c;
8'h85 : rvCrc[2] <= 32'heaec5d1b;
8'h86 : rvCrc[2] <= 32'he885a892;
8'h87 : rvCrc[2] <= 32'he95d0415;
8'h88 : rvCrc[2] <= 32'he29327b8;
8'h89 : rvCrc[2] <= 32'he34b8b3f;
8'h8a : rvCrc[2] <= 32'he1227eb6;
8'h8b : rvCrc[2] <= 32'he0fad231;
8'h8c : rvCrc[2] <= 32'he5f195a4;
8'h8d : rvCrc[2] <= 32'he4293923;
8'h8e : rvCrc[2] <= 32'he640ccaa;
8'h8f : rvCrc[2] <= 32'he798602d;
8'h90 : rvCrc[2] <= 32'hf1dc8bf0;
8'h91 : rvCrc[2] <= 32'hf0042777;
8'h92 : rvCrc[2] <= 32'hf26dd2fe;
8'h93 : rvCrc[2] <= 32'hf3b57e79;
8'h94 : rvCrc[2] <= 32'hf6be39ec;
8'h95 : rvCrc[2] <= 32'hf766956b;
8'h96 : rvCrc[2] <= 32'hf50f60e2;
8'h97 : rvCrc[2] <= 32'hf4d7cc65;
8'h98 : rvCrc[2] <= 32'hff19efc8;
8'h99 : rvCrc[2] <= 32'hfec1434f;
8'h9a : rvCrc[2] <= 32'hfca8b6c6;
8'h9b : rvCrc[2] <= 32'hfd701a41;
8'h9c : rvCrc[2] <= 32'hf87b5dd4;
8'h9d : rvCrc[2] <= 32'hf9a3f153;
8'h9e : rvCrc[2] <= 32'hfbca04da;
8'h9f : rvCrc[2] <= 32'hfa12a85d;
8'ha0 : rvCrc[2] <= 32'hd743d360;
8'ha1 : rvCrc[2] <= 32'hd69b7fe7;
8'ha2 : rvCrc[2] <= 32'hd4f28a6e;
8'ha3 : rvCrc[2] <= 32'hd52a26e9;
8'ha4 : rvCrc[2] <= 32'hd021617c;
8'ha5 : rvCrc[2] <= 32'hd1f9cdfb;
8'ha6 : rvCrc[2] <= 32'hd3903872;
8'ha7 : rvCrc[2] <= 32'hd24894f5;
8'ha8 : rvCrc[2] <= 32'hd986b758;
8'ha9 : rvCrc[2] <= 32'hd85e1bdf;
8'haa : rvCrc[2] <= 32'hda37ee56;
8'hab : rvCrc[2] <= 32'hdbef42d1;
8'hac : rvCrc[2] <= 32'hdee40544;
8'had : rvCrc[2] <= 32'hdf3ca9c3;
8'hae : rvCrc[2] <= 32'hdd555c4a;
8'haf : rvCrc[2] <= 32'hdc8df0cd;
8'hb0 : rvCrc[2] <= 32'hcac91b10;
8'hb1 : rvCrc[2] <= 32'hcb11b797;
8'hb2 : rvCrc[2] <= 32'hc978421e;
8'hb3 : rvCrc[2] <= 32'hc8a0ee99;
8'hb4 : rvCrc[2] <= 32'hcdaba90c;
8'hb5 : rvCrc[2] <= 32'hcc73058b;
8'hb6 : rvCrc[2] <= 32'hce1af002;
8'hb7 : rvCrc[2] <= 32'hcfc25c85;
8'hb8 : rvCrc[2] <= 32'hc40c7f28;
8'hb9 : rvCrc[2] <= 32'hc5d4d3af;
8'hba : rvCrc[2] <= 32'hc7bd2626;
8'hbb : rvCrc[2] <= 32'hc6658aa1;
8'hbc : rvCrc[2] <= 32'hc36ecd34;
8'hbd : rvCrc[2] <= 32'hc2b661b3;
8'hbe : rvCrc[2] <= 32'hc0df943a;
8'hbf : rvCrc[2] <= 32'hc10738bd;
8'hc0 : rvCrc[2] <= 32'h9a7d6240;
8'hc1 : rvCrc[2] <= 32'h9ba5cec7;
8'hc2 : rvCrc[2] <= 32'h99cc3b4e;
8'hc3 : rvCrc[2] <= 32'h981497c9;
8'hc4 : rvCrc[2] <= 32'h9d1fd05c;
8'hc5 : rvCrc[2] <= 32'h9cc77cdb;
8'hc6 : rvCrc[2] <= 32'h9eae8952;
8'hc7 : rvCrc[2] <= 32'h9f7625d5;
8'hc8 : rvCrc[2] <= 32'h94b80678;
8'hc9 : rvCrc[2] <= 32'h9560aaff;
8'hca : rvCrc[2] <= 32'h97095f76;
8'hcb : rvCrc[2] <= 32'h96d1f3f1;
8'hcc : rvCrc[2] <= 32'h93dab464;
8'hcd : rvCrc[2] <= 32'h920218e3;
8'hce : rvCrc[2] <= 32'h906bed6a;
8'hcf : rvCrc[2] <= 32'h91b341ed;
8'hd0 : rvCrc[2] <= 32'h87f7aa30;
8'hd1 : rvCrc[2] <= 32'h862f06b7;
8'hd2 : rvCrc[2] <= 32'h8446f33e;
8'hd3 : rvCrc[2] <= 32'h859e5fb9;
8'hd4 : rvCrc[2] <= 32'h8095182c;
8'hd5 : rvCrc[2] <= 32'h814db4ab;
8'hd6 : rvCrc[2] <= 32'h83244122;
8'hd7 : rvCrc[2] <= 32'h82fceda5;
8'hd8 : rvCrc[2] <= 32'h8932ce08;
8'hd9 : rvCrc[2] <= 32'h88ea628f;
8'hda : rvCrc[2] <= 32'h8a839706;
8'hdb : rvCrc[2] <= 32'h8b5b3b81;
8'hdc : rvCrc[2] <= 32'h8e507c14;
8'hdd : rvCrc[2] <= 32'h8f88d093;
8'hde : rvCrc[2] <= 32'h8de1251a;
8'hdf : rvCrc[2] <= 32'h8c39899d;
8'he0 : rvCrc[2] <= 32'ha168f2a0;
8'he1 : rvCrc[2] <= 32'ha0b05e27;
8'he2 : rvCrc[2] <= 32'ha2d9abae;
8'he3 : rvCrc[2] <= 32'ha3010729;
8'he4 : rvCrc[2] <= 32'ha60a40bc;
8'he5 : rvCrc[2] <= 32'ha7d2ec3b;
8'he6 : rvCrc[2] <= 32'ha5bb19b2;
8'he7 : rvCrc[2] <= 32'ha463b535;
8'he8 : rvCrc[2] <= 32'hafad9698;
8'he9 : rvCrc[2] <= 32'hae753a1f;
8'hea : rvCrc[2] <= 32'hac1ccf96;
8'heb : rvCrc[2] <= 32'hadc46311;
8'hec : rvCrc[2] <= 32'ha8cf2484;
8'hed : rvCrc[2] <= 32'ha9178803;
8'hee : rvCrc[2] <= 32'hab7e7d8a;
8'hef : rvCrc[2] <= 32'haaa6d10d;
8'hf0 : rvCrc[2] <= 32'hbce23ad0;
8'hf1 : rvCrc[2] <= 32'hbd3a9657;
8'hf2 : rvCrc[2] <= 32'hbf5363de;
8'hf3 : rvCrc[2] <= 32'hbe8bcf59;
8'hf4 : rvCrc[2] <= 32'hbb8088cc;
8'hf5 : rvCrc[2] <= 32'hba58244b;
8'hf6 : rvCrc[2] <= 32'hb831d1c2;
8'hf7 : rvCrc[2] <= 32'hb9e97d45;
8'hf8 : rvCrc[2] <= 32'hb2275ee8;
8'hf9 : rvCrc[2] <= 32'hb3fff26f;
8'hfa : rvCrc[2] <= 32'hb19607e6;
8'hfb : rvCrc[2] <= 32'hb04eab61;
8'hfc : rvCrc[2] <= 32'hb545ecf4;
8'hfd : rvCrc[2] <= 32'hb49d4073;
8'hfe : rvCrc[2] <= 32'hb6f4b5fa;
8'hff : rvCrc[2] <= 32'hb72c197d;
endcase
case(iv_Input[031:024])
8'h00 : rvCrc[3] <= 32'h00000000;
8'h01 : rvCrc[3] <= 32'hdc6d9ab7;
8'h02 : rvCrc[3] <= 32'hbc1a28d9;
8'h03 : rvCrc[3] <= 32'h6077b26e;
8'h04 : rvCrc[3] <= 32'h7cf54c05;
8'h05 : rvCrc[3] <= 32'ha098d6b2;
8'h06 : rvCrc[3] <= 32'hc0ef64dc;
8'h07 : rvCrc[3] <= 32'h1c82fe6b;
8'h08 : rvCrc[3] <= 32'hf9ea980a;
8'h09 : rvCrc[3] <= 32'h258702bd;
8'h0a : rvCrc[3] <= 32'h45f0b0d3;
8'h0b : rvCrc[3] <= 32'h999d2a64;
8'h0c : rvCrc[3] <= 32'h851fd40f;
8'h0d : rvCrc[3] <= 32'h59724eb8;
8'h0e : rvCrc[3] <= 32'h3905fcd6;
8'h0f : rvCrc[3] <= 32'he5686661;
8'h10 : rvCrc[3] <= 32'hf7142da3;
8'h11 : rvCrc[3] <= 32'h2b79b714;
8'h12 : rvCrc[3] <= 32'h4b0e057a;
8'h13 : rvCrc[3] <= 32'h97639fcd;
8'h14 : rvCrc[3] <= 32'h8be161a6;
8'h15 : rvCrc[3] <= 32'h578cfb11;
8'h16 : rvCrc[3] <= 32'h37fb497f;
8'h17 : rvCrc[3] <= 32'heb96d3c8;
8'h18 : rvCrc[3] <= 32'h0efeb5a9;
8'h19 : rvCrc[3] <= 32'hd2932f1e;
8'h1a : rvCrc[3] <= 32'hb2e49d70;
8'h1b : rvCrc[3] <= 32'h6e8907c7;
8'h1c : rvCrc[3] <= 32'h720bf9ac;
8'h1d : rvCrc[3] <= 32'hae66631b;
8'h1e : rvCrc[3] <= 32'hce11d175;
8'h1f : rvCrc[3] <= 32'h127c4bc2;
8'h20 : rvCrc[3] <= 32'heae946f1;
8'h21 : rvCrc[3] <= 32'h3684dc46;
8'h22 : rvCrc[3] <= 32'h56f36e28;
8'h23 : rvCrc[3] <= 32'h8a9ef49f;
8'h24 : rvCrc[3] <= 32'h961c0af4;
8'h25 : rvCrc[3] <= 32'h4a719043;
8'h26 : rvCrc[3] <= 32'h2a06222d;
8'h27 : rvCrc[3] <= 32'hf66bb89a;
8'h28 : rvCrc[3] <= 32'h1303defb;
8'h29 : rvCrc[3] <= 32'hcf6e444c;
8'h2a : rvCrc[3] <= 32'haf19f622;
8'h2b : rvCrc[3] <= 32'h73746c95;
8'h2c : rvCrc[3] <= 32'h6ff692fe;
8'h2d : rvCrc[3] <= 32'hb39b0849;
8'h2e : rvCrc[3] <= 32'hd3ecba27;
8'h2f : rvCrc[3] <= 32'h0f812090;
8'h30 : rvCrc[3] <= 32'h1dfd6b52;
8'h31 : rvCrc[3] <= 32'hc190f1e5;
8'h32 : rvCrc[3] <= 32'ha1e7438b;
8'h33 : rvCrc[3] <= 32'h7d8ad93c;
8'h34 : rvCrc[3] <= 32'h61082757;
8'h35 : rvCrc[3] <= 32'hbd65bde0;
8'h36 : rvCrc[3] <= 32'hdd120f8e;
8'h37 : rvCrc[3] <= 32'h017f9539;
8'h38 : rvCrc[3] <= 32'he417f358;
8'h39 : rvCrc[3] <= 32'h387a69ef;
8'h3a : rvCrc[3] <= 32'h580ddb81;
8'h3b : rvCrc[3] <= 32'h84604136;
8'h3c : rvCrc[3] <= 32'h98e2bf5d;
8'h3d : rvCrc[3] <= 32'h448f25ea;
8'h3e : rvCrc[3] <= 32'h24f89784;
8'h3f : rvCrc[3] <= 32'hf8950d33;
8'h40 : rvCrc[3] <= 32'hd1139055;
8'h41 : rvCrc[3] <= 32'h0d7e0ae2;
8'h42 : rvCrc[3] <= 32'h6d09b88c;
8'h43 : rvCrc[3] <= 32'hb164223b;
8'h44 : rvCrc[3] <= 32'hade6dc50;
8'h45 : rvCrc[3] <= 32'h718b46e7;
8'h46 : rvCrc[3] <= 32'h11fcf489;
8'h47 : rvCrc[3] <= 32'hcd916e3e;
8'h48 : rvCrc[3] <= 32'h28f9085f;
8'h49 : rvCrc[3] <= 32'hf49492e8;
8'h4a : rvCrc[3] <= 32'h94e32086;
8'h4b : rvCrc[3] <= 32'h488eba31;
8'h4c : rvCrc[3] <= 32'h540c445a;
8'h4d : rvCrc[3] <= 32'h8861deed;
8'h4e : rvCrc[3] <= 32'he8166c83;
8'h4f : rvCrc[3] <= 32'h347bf634;
8'h50 : rvCrc[3] <= 32'h2607bdf6;
8'h51 : rvCrc[3] <= 32'hfa6a2741;
8'h52 : rvCrc[3] <= 32'h9a1d952f;
8'h53 : rvCrc[3] <= 32'h46700f98;
8'h54 : rvCrc[3] <= 32'h5af2f1f3;
8'h55 : rvCrc[3] <= 32'h869f6b44;
8'h56 : rvCrc[3] <= 32'he6e8d92a;
8'h57 : rvCrc[3] <= 32'h3a85439d;
8'h58 : rvCrc[3] <= 32'hdfed25fc;
8'h59 : rvCrc[3] <= 32'h0380bf4b;
8'h5a : rvCrc[3] <= 32'h63f70d25;
8'h5b : rvCrc[3] <= 32'hbf9a9792;
8'h5c : rvCrc[3] <= 32'ha31869f9;
8'h5d : rvCrc[3] <= 32'h7f75f34e;
8'h5e : rvCrc[3] <= 32'h1f024120;
8'h5f : rvCrc[3] <= 32'hc36fdb97;
8'h60 : rvCrc[3] <= 32'h3bfad6a4;
8'h61 : rvCrc[3] <= 32'he7974c13;
8'h62 : rvCrc[3] <= 32'h87e0fe7d;
8'h63 : rvCrc[3] <= 32'h5b8d64ca;
8'h64 : rvCrc[3] <= 32'h470f9aa1;
8'h65 : rvCrc[3] <= 32'h9b620016;
8'h66 : rvCrc[3] <= 32'hfb15b278;
8'h67 : rvCrc[3] <= 32'h277828cf;
8'h68 : rvCrc[3] <= 32'hc2104eae;
8'h69 : rvCrc[3] <= 32'h1e7dd419;
8'h6a : rvCrc[3] <= 32'h7e0a6677;
8'h6b : rvCrc[3] <= 32'ha267fcc0;
8'h6c : rvCrc[3] <= 32'hbee502ab;
8'h6d : rvCrc[3] <= 32'h6288981c;
8'h6e : rvCrc[3] <= 32'h02ff2a72;
8'h6f : rvCrc[3] <= 32'hde92b0c5;
8'h70 : rvCrc[3] <= 32'hcceefb07;
8'h71 : rvCrc[3] <= 32'h108361b0;
8'h72 : rvCrc[3] <= 32'h70f4d3de;
8'h73 : rvCrc[3] <= 32'hac994969;
8'h74 : rvCrc[3] <= 32'hb01bb702;
8'h75 : rvCrc[3] <= 32'h6c762db5;
8'h76 : rvCrc[3] <= 32'h0c019fdb;
8'h77 : rvCrc[3] <= 32'hd06c056c;
8'h78 : rvCrc[3] <= 32'h3504630d;
8'h79 : rvCrc[3] <= 32'he969f9ba;
8'h7a : rvCrc[3] <= 32'h891e4bd4;
8'h7b : rvCrc[3] <= 32'h5573d163;
8'h7c : rvCrc[3] <= 32'h49f12f08;
8'h7d : rvCrc[3] <= 32'h959cb5bf;
8'h7e : rvCrc[3] <= 32'hf5eb07d1;
8'h7f : rvCrc[3] <= 32'h29869d66;
8'h80 : rvCrc[3] <= 32'ha6e63d1d;
8'h81 : rvCrc[3] <= 32'h7a8ba7aa;
8'h82 : rvCrc[3] <= 32'h1afc15c4;
8'h83 : rvCrc[3] <= 32'hc6918f73;
8'h84 : rvCrc[3] <= 32'hda137118;
8'h85 : rvCrc[3] <= 32'h067eebaf;
8'h86 : rvCrc[3] <= 32'h660959c1;
8'h87 : rvCrc[3] <= 32'hba64c376;
8'h88 : rvCrc[3] <= 32'h5f0ca517;
8'h89 : rvCrc[3] <= 32'h83613fa0;
8'h8a : rvCrc[3] <= 32'he3168dce;
8'h8b : rvCrc[3] <= 32'h3f7b1779;
8'h8c : rvCrc[3] <= 32'h23f9e912;
8'h8d : rvCrc[3] <= 32'hff9473a5;
8'h8e : rvCrc[3] <= 32'h9fe3c1cb;
8'h8f : rvCrc[3] <= 32'h438e5b7c;
8'h90 : rvCrc[3] <= 32'h51f210be;
8'h91 : rvCrc[3] <= 32'h8d9f8a09;
8'h92 : rvCrc[3] <= 32'hede83867;
8'h93 : rvCrc[3] <= 32'h3185a2d0;
8'h94 : rvCrc[3] <= 32'h2d075cbb;
8'h95 : rvCrc[3] <= 32'hf16ac60c;
8'h96 : rvCrc[3] <= 32'h911d7462;
8'h97 : rvCrc[3] <= 32'h4d70eed5;
8'h98 : rvCrc[3] <= 32'ha81888b4;
8'h99 : rvCrc[3] <= 32'h74751203;
8'h9a : rvCrc[3] <= 32'h1402a06d;
8'h9b : rvCrc[3] <= 32'hc86f3ada;
8'h9c : rvCrc[3] <= 32'hd4edc4b1;
8'h9d : rvCrc[3] <= 32'h08805e06;
8'h9e : rvCrc[3] <= 32'h68f7ec68;
8'h9f : rvCrc[3] <= 32'hb49a76df;
8'ha0 : rvCrc[3] <= 32'h4c0f7bec;
8'ha1 : rvCrc[3] <= 32'h9062e15b;
8'ha2 : rvCrc[3] <= 32'hf0155335;
8'ha3 : rvCrc[3] <= 32'h2c78c982;
8'ha4 : rvCrc[3] <= 32'h30fa37e9;
8'ha5 : rvCrc[3] <= 32'hec97ad5e;
8'ha6 : rvCrc[3] <= 32'h8ce01f30;
8'ha7 : rvCrc[3] <= 32'h508d8587;
8'ha8 : rvCrc[3] <= 32'hb5e5e3e6;
8'ha9 : rvCrc[3] <= 32'h69887951;
8'haa : rvCrc[3] <= 32'h09ffcb3f;
8'hab : rvCrc[3] <= 32'hd5925188;
8'hac : rvCrc[3] <= 32'hc910afe3;
8'had : rvCrc[3] <= 32'h157d3554;
8'hae : rvCrc[3] <= 32'h750a873a;
8'haf : rvCrc[3] <= 32'ha9671d8d;
8'hb0 : rvCrc[3] <= 32'hbb1b564f;
8'hb1 : rvCrc[3] <= 32'h6776ccf8;
8'hb2 : rvCrc[3] <= 32'h07017e96;
8'hb3 : rvCrc[3] <= 32'hdb6ce421;
8'hb4 : rvCrc[3] <= 32'hc7ee1a4a;
8'hb5 : rvCrc[3] <= 32'h1b8380fd;
8'hb6 : rvCrc[3] <= 32'h7bf43293;
8'hb7 : rvCrc[3] <= 32'ha799a824;
8'hb8 : rvCrc[3] <= 32'h42f1ce45;
8'hb9 : rvCrc[3] <= 32'h9e9c54f2;
8'hba : rvCrc[3] <= 32'hfeebe69c;
8'hbb : rvCrc[3] <= 32'h22867c2b;
8'hbc : rvCrc[3] <= 32'h3e048240;
8'hbd : rvCrc[3] <= 32'he26918f7;
8'hbe : rvCrc[3] <= 32'h821eaa99;
8'hbf : rvCrc[3] <= 32'h5e73302e;
8'hc0 : rvCrc[3] <= 32'h77f5ad48;
8'hc1 : rvCrc[3] <= 32'hab9837ff;
8'hc2 : rvCrc[3] <= 32'hcbef8591;
8'hc3 : rvCrc[3] <= 32'h17821f26;
8'hc4 : rvCrc[3] <= 32'h0b00e14d;
8'hc5 : rvCrc[3] <= 32'hd76d7bfa;
8'hc6 : rvCrc[3] <= 32'hb71ac994;
8'hc7 : rvCrc[3] <= 32'h6b775323;
8'hc8 : rvCrc[3] <= 32'h8e1f3542;
8'hc9 : rvCrc[3] <= 32'h5272aff5;
8'hca : rvCrc[3] <= 32'h32051d9b;
8'hcb : rvCrc[3] <= 32'hee68872c;
8'hcc : rvCrc[3] <= 32'hf2ea7947;
8'hcd : rvCrc[3] <= 32'h2e87e3f0;
8'hce : rvCrc[3] <= 32'h4ef0519e;
8'hcf : rvCrc[3] <= 32'h929dcb29;
8'hd0 : rvCrc[3] <= 32'h80e180eb;
8'hd1 : rvCrc[3] <= 32'h5c8c1a5c;
8'hd2 : rvCrc[3] <= 32'h3cfba832;
8'hd3 : rvCrc[3] <= 32'he0963285;
8'hd4 : rvCrc[3] <= 32'hfc14ccee;
8'hd5 : rvCrc[3] <= 32'h20795659;
8'hd6 : rvCrc[3] <= 32'h400ee437;
8'hd7 : rvCrc[3] <= 32'h9c637e80;
8'hd8 : rvCrc[3] <= 32'h790b18e1;
8'hd9 : rvCrc[3] <= 32'ha5668256;
8'hda : rvCrc[3] <= 32'hc5113038;
8'hdb : rvCrc[3] <= 32'h197caa8f;
8'hdc : rvCrc[3] <= 32'h05fe54e4;
8'hdd : rvCrc[3] <= 32'hd993ce53;
8'hde : rvCrc[3] <= 32'hb9e47c3d;
8'hdf : rvCrc[3] <= 32'h6589e68a;
8'he0 : rvCrc[3] <= 32'h9d1cebb9;
8'he1 : rvCrc[3] <= 32'h4171710e;
8'he2 : rvCrc[3] <= 32'h2106c360;
8'he3 : rvCrc[3] <= 32'hfd6b59d7;
8'he4 : rvCrc[3] <= 32'he1e9a7bc;
8'he5 : rvCrc[3] <= 32'h3d843d0b;
8'he6 : rvCrc[3] <= 32'h5df38f65;
8'he7 : rvCrc[3] <= 32'h819e15d2;
8'he8 : rvCrc[3] <= 32'h64f673b3;
8'he9 : rvCrc[3] <= 32'hb89be904;
8'hea : rvCrc[3] <= 32'hd8ec5b6a;
8'heb : rvCrc[3] <= 32'h0481c1dd;
8'hec : rvCrc[3] <= 32'h18033fb6;
8'hed : rvCrc[3] <= 32'hc46ea501;
8'hee : rvCrc[3] <= 32'ha419176f;
8'hef : rvCrc[3] <= 32'h78748dd8;
8'hf0 : rvCrc[3] <= 32'h6a08c61a;
8'hf1 : rvCrc[3] <= 32'hb6655cad;
8'hf2 : rvCrc[3] <= 32'hd612eec3;
8'hf3 : rvCrc[3] <= 32'h0a7f7474;
8'hf4 : rvCrc[3] <= 32'h16fd8a1f;
8'hf5 : rvCrc[3] <= 32'hca9010a8;
8'hf6 : rvCrc[3] <= 32'haae7a2c6;
8'hf7 : rvCrc[3] <= 32'h768a3871;
8'hf8 : rvCrc[3] <= 32'h93e25e10;
8'hf9 : rvCrc[3] <= 32'h4f8fc4a7;
8'hfa : rvCrc[3] <= 32'h2ff876c9;
8'hfb : rvCrc[3] <= 32'hf395ec7e;
8'hfc : rvCrc[3] <= 32'hef171215;
8'hfd : rvCrc[3] <= 32'h337a88a2;
8'hfe : rvCrc[3] <= 32'h530d3acc;
8'hff : rvCrc[3] <= 32'h8f60a07b;
endcase
case(iv_Input[039:032])
8'h00 : rvCrc[4] <= 32'h00000000;
8'h01 : rvCrc[4] <= 32'h490d678d;
8'h02 : rvCrc[4] <= 32'h921acf1a;
8'h03 : rvCrc[4] <= 32'hdb17a897;
8'h04 : rvCrc[4] <= 32'h20f48383;
8'h05 : rvCrc[4] <= 32'h69f9e40e;
8'h06 : rvCrc[4] <= 32'hb2ee4c99;
8'h07 : rvCrc[4] <= 32'hfbe32b14;
8'h08 : rvCrc[4] <= 32'h41e90706;
8'h09 : rvCrc[4] <= 32'h08e4608b;
8'h0a : rvCrc[4] <= 32'hd3f3c81c;
8'h0b : rvCrc[4] <= 32'h9afeaf91;
8'h0c : rvCrc[4] <= 32'h611d8485;
8'h0d : rvCrc[4] <= 32'h2810e308;
8'h0e : rvCrc[4] <= 32'hf3074b9f;
8'h0f : rvCrc[4] <= 32'hba0a2c12;
8'h10 : rvCrc[4] <= 32'h83d20e0c;
8'h11 : rvCrc[4] <= 32'hcadf6981;
8'h12 : rvCrc[4] <= 32'h11c8c116;
8'h13 : rvCrc[4] <= 32'h58c5a69b;
8'h14 : rvCrc[4] <= 32'ha3268d8f;
8'h15 : rvCrc[4] <= 32'hea2bea02;
8'h16 : rvCrc[4] <= 32'h313c4295;
8'h17 : rvCrc[4] <= 32'h78312518;
8'h18 : rvCrc[4] <= 32'hc23b090a;
8'h19 : rvCrc[4] <= 32'h8b366e87;
8'h1a : rvCrc[4] <= 32'h5021c610;
8'h1b : rvCrc[4] <= 32'h192ca19d;
8'h1c : rvCrc[4] <= 32'he2cf8a89;
8'h1d : rvCrc[4] <= 32'habc2ed04;
8'h1e : rvCrc[4] <= 32'h70d54593;
8'h1f : rvCrc[4] <= 32'h39d8221e;
8'h20 : rvCrc[4] <= 32'h036501af;
8'h21 : rvCrc[4] <= 32'h4a686622;
8'h22 : rvCrc[4] <= 32'h917fceb5;
8'h23 : rvCrc[4] <= 32'hd872a938;
8'h24 : rvCrc[4] <= 32'h2391822c;
8'h25 : rvCrc[4] <= 32'h6a9ce5a1;
8'h26 : rvCrc[4] <= 32'hb18b4d36;
8'h27 : rvCrc[4] <= 32'hf8862abb;
8'h28 : rvCrc[4] <= 32'h428c06a9;
8'h29 : rvCrc[4] <= 32'h0b816124;
8'h2a : rvCrc[4] <= 32'hd096c9b3;
8'h2b : rvCrc[4] <= 32'h999bae3e;
8'h2c : rvCrc[4] <= 32'h6278852a;
8'h2d : rvCrc[4] <= 32'h2b75e2a7;
8'h2e : rvCrc[4] <= 32'hf0624a30;
8'h2f : rvCrc[4] <= 32'hb96f2dbd;
8'h30 : rvCrc[4] <= 32'h80b70fa3;
8'h31 : rvCrc[4] <= 32'hc9ba682e;
8'h32 : rvCrc[4] <= 32'h12adc0b9;
8'h33 : rvCrc[4] <= 32'h5ba0a734;
8'h34 : rvCrc[4] <= 32'ha0438c20;
8'h35 : rvCrc[4] <= 32'he94eebad;
8'h36 : rvCrc[4] <= 32'h3259433a;
8'h37 : rvCrc[4] <= 32'h7b5424b7;
8'h38 : rvCrc[4] <= 32'hc15e08a5;
8'h39 : rvCrc[4] <= 32'h88536f28;
8'h3a : rvCrc[4] <= 32'h5344c7bf;
8'h3b : rvCrc[4] <= 32'h1a49a032;
8'h3c : rvCrc[4] <= 32'he1aa8b26;
8'h3d : rvCrc[4] <= 32'ha8a7ecab;
8'h3e : rvCrc[4] <= 32'h73b0443c;
8'h3f : rvCrc[4] <= 32'h3abd23b1;
8'h40 : rvCrc[4] <= 32'h06ca035e;
8'h41 : rvCrc[4] <= 32'h4fc764d3;
8'h42 : rvCrc[4] <= 32'h94d0cc44;
8'h43 : rvCrc[4] <= 32'hddddabc9;
8'h44 : rvCrc[4] <= 32'h263e80dd;
8'h45 : rvCrc[4] <= 32'h6f33e750;
8'h46 : rvCrc[4] <= 32'hb4244fc7;
8'h47 : rvCrc[4] <= 32'hfd29284a;
8'h48 : rvCrc[4] <= 32'h47230458;
8'h49 : rvCrc[4] <= 32'h0e2e63d5;
8'h4a : rvCrc[4] <= 32'hd539cb42;
8'h4b : rvCrc[4] <= 32'h9c34accf;
8'h4c : rvCrc[4] <= 32'h67d787db;
8'h4d : rvCrc[4] <= 32'h2edae056;
8'h4e : rvCrc[4] <= 32'hf5cd48c1;
8'h4f : rvCrc[4] <= 32'hbcc02f4c;
8'h50 : rvCrc[4] <= 32'h85180d52;
8'h51 : rvCrc[4] <= 32'hcc156adf;
8'h52 : rvCrc[4] <= 32'h1702c248;
8'h53 : rvCrc[4] <= 32'h5e0fa5c5;
8'h54 : rvCrc[4] <= 32'ha5ec8ed1;
8'h55 : rvCrc[4] <= 32'hece1e95c;
8'h56 : rvCrc[4] <= 32'h37f641cb;
8'h57 : rvCrc[4] <= 32'h7efb2646;
8'h58 : rvCrc[4] <= 32'hc4f10a54;
8'h59 : rvCrc[4] <= 32'h8dfc6dd9;
8'h5a : rvCrc[4] <= 32'h56ebc54e;
8'h5b : rvCrc[4] <= 32'h1fe6a2c3;
8'h5c : rvCrc[4] <= 32'he40589d7;
8'h5d : rvCrc[4] <= 32'had08ee5a;
8'h5e : rvCrc[4] <= 32'h761f46cd;
8'h5f : rvCrc[4] <= 32'h3f122140;
8'h60 : rvCrc[4] <= 32'h05af02f1;
8'h61 : rvCrc[4] <= 32'h4ca2657c;
8'h62 : rvCrc[4] <= 32'h97b5cdeb;
8'h63 : rvCrc[4] <= 32'hdeb8aa66;
8'h64 : rvCrc[4] <= 32'h255b8172;
8'h65 : rvCrc[4] <= 32'h6c56e6ff;
8'h66 : rvCrc[4] <= 32'hb7414e68;
8'h67 : rvCrc[4] <= 32'hfe4c29e5;
8'h68 : rvCrc[4] <= 32'h444605f7;
8'h69 : rvCrc[4] <= 32'h0d4b627a;
8'h6a : rvCrc[4] <= 32'hd65ccaed;
8'h6b : rvCrc[4] <= 32'h9f51ad60;
8'h6c : rvCrc[4] <= 32'h64b28674;
8'h6d : rvCrc[4] <= 32'h2dbfe1f9;
8'h6e : rvCrc[4] <= 32'hf6a8496e;
8'h6f : rvCrc[4] <= 32'hbfa52ee3;
8'h70 : rvCrc[4] <= 32'h867d0cfd;
8'h71 : rvCrc[4] <= 32'hcf706b70;
8'h72 : rvCrc[4] <= 32'h1467c3e7;
8'h73 : rvCrc[4] <= 32'h5d6aa46a;
8'h74 : rvCrc[4] <= 32'ha6898f7e;
8'h75 : rvCrc[4] <= 32'hef84e8f3;
8'h76 : rvCrc[4] <= 32'h34934064;
8'h77 : rvCrc[4] <= 32'h7d9e27e9;
8'h78 : rvCrc[4] <= 32'hc7940bfb;
8'h79 : rvCrc[4] <= 32'h8e996c76;
8'h7a : rvCrc[4] <= 32'h558ec4e1;
8'h7b : rvCrc[4] <= 32'h1c83a36c;
8'h7c : rvCrc[4] <= 32'he7608878;
8'h7d : rvCrc[4] <= 32'hae6deff5;
8'h7e : rvCrc[4] <= 32'h757a4762;
8'h7f : rvCrc[4] <= 32'h3c7720ef;
8'h80 : rvCrc[4] <= 32'h0d9406bc;
8'h81 : rvCrc[4] <= 32'h44996131;
8'h82 : rvCrc[4] <= 32'h9f8ec9a6;
8'h83 : rvCrc[4] <= 32'hd683ae2b;
8'h84 : rvCrc[4] <= 32'h2d60853f;
8'h85 : rvCrc[4] <= 32'h646de2b2;
8'h86 : rvCrc[4] <= 32'hbf7a4a25;
8'h87 : rvCrc[4] <= 32'hf6772da8;
8'h88 : rvCrc[4] <= 32'h4c7d01ba;
8'h89 : rvCrc[4] <= 32'h05706637;
8'h8a : rvCrc[4] <= 32'hde67cea0;
8'h8b : rvCrc[4] <= 32'h976aa92d;
8'h8c : rvCrc[4] <= 32'h6c898239;
8'h8d : rvCrc[4] <= 32'h2584e5b4;
8'h8e : rvCrc[4] <= 32'hfe934d23;
8'h8f : rvCrc[4] <= 32'hb79e2aae;
8'h90 : rvCrc[4] <= 32'h8e4608b0;
8'h91 : rvCrc[4] <= 32'hc74b6f3d;
8'h92 : rvCrc[4] <= 32'h1c5cc7aa;
8'h93 : rvCrc[4] <= 32'h5551a027;
8'h94 : rvCrc[4] <= 32'haeb28b33;
8'h95 : rvCrc[4] <= 32'he7bfecbe;
8'h96 : rvCrc[4] <= 32'h3ca84429;
8'h97 : rvCrc[4] <= 32'h75a523a4;
8'h98 : rvCrc[4] <= 32'hcfaf0fb6;
8'h99 : rvCrc[4] <= 32'h86a2683b;
8'h9a : rvCrc[4] <= 32'h5db5c0ac;
8'h9b : rvCrc[4] <= 32'h14b8a721;
8'h9c : rvCrc[4] <= 32'hef5b8c35;
8'h9d : rvCrc[4] <= 32'ha656ebb8;
8'h9e : rvCrc[4] <= 32'h7d41432f;
8'h9f : rvCrc[4] <= 32'h344c24a2;
8'ha0 : rvCrc[4] <= 32'h0ef10713;
8'ha1 : rvCrc[4] <= 32'h47fc609e;
8'ha2 : rvCrc[4] <= 32'h9cebc809;
8'ha3 : rvCrc[4] <= 32'hd5e6af84;
8'ha4 : rvCrc[4] <= 32'h2e058490;
8'ha5 : rvCrc[4] <= 32'h6708e31d;
8'ha6 : rvCrc[4] <= 32'hbc1f4b8a;
8'ha7 : rvCrc[4] <= 32'hf5122c07;
8'ha8 : rvCrc[4] <= 32'h4f180015;
8'ha9 : rvCrc[4] <= 32'h06156798;
8'haa : rvCrc[4] <= 32'hdd02cf0f;
8'hab : rvCrc[4] <= 32'h940fa882;
8'hac : rvCrc[4] <= 32'h6fec8396;
8'had : rvCrc[4] <= 32'h26e1e41b;
8'hae : rvCrc[4] <= 32'hfdf64c8c;
8'haf : rvCrc[4] <= 32'hb4fb2b01;
8'hb0 : rvCrc[4] <= 32'h8d23091f;
8'hb1 : rvCrc[4] <= 32'hc42e6e92;
8'hb2 : rvCrc[4] <= 32'h1f39c605;
8'hb3 : rvCrc[4] <= 32'h5634a188;
8'hb4 : rvCrc[4] <= 32'hadd78a9c;
8'hb5 : rvCrc[4] <= 32'he4daed11;
8'hb6 : rvCrc[4] <= 32'h3fcd4586;
8'hb7 : rvCrc[4] <= 32'h76c0220b;
8'hb8 : rvCrc[4] <= 32'hccca0e19;
8'hb9 : rvCrc[4] <= 32'h85c76994;
8'hba : rvCrc[4] <= 32'h5ed0c103;
8'hbb : rvCrc[4] <= 32'h17dda68e;
8'hbc : rvCrc[4] <= 32'hec3e8d9a;
8'hbd : rvCrc[4] <= 32'ha533ea17;
8'hbe : rvCrc[4] <= 32'h7e244280;
8'hbf : rvCrc[4] <= 32'h3729250d;
8'hc0 : rvCrc[4] <= 32'h0b5e05e2;
8'hc1 : rvCrc[4] <= 32'h4253626f;
8'hc2 : rvCrc[4] <= 32'h9944caf8;
8'hc3 : rvCrc[4] <= 32'hd049ad75;
8'hc4 : rvCrc[4] <= 32'h2baa8661;
8'hc5 : rvCrc[4] <= 32'h62a7e1ec;
8'hc6 : rvCrc[4] <= 32'hb9b0497b;
8'hc7 : rvCrc[4] <= 32'hf0bd2ef6;
8'hc8 : rvCrc[4] <= 32'h4ab702e4;
8'hc9 : rvCrc[4] <= 32'h03ba6569;
8'hca : rvCrc[4] <= 32'hd8adcdfe;
8'hcb : rvCrc[4] <= 32'h91a0aa73;
8'hcc : rvCrc[4] <= 32'h6a438167;
8'hcd : rvCrc[4] <= 32'h234ee6ea;
8'hce : rvCrc[4] <= 32'hf8594e7d;
8'hcf : rvCrc[4] <= 32'hb15429f0;
8'hd0 : rvCrc[4] <= 32'h888c0bee;
8'hd1 : rvCrc[4] <= 32'hc1816c63;
8'hd2 : rvCrc[4] <= 32'h1a96c4f4;
8'hd3 : rvCrc[4] <= 32'h539ba379;
8'hd4 : rvCrc[4] <= 32'ha878886d;
8'hd5 : rvCrc[4] <= 32'he175efe0;
8'hd6 : rvCrc[4] <= 32'h3a624777;
8'hd7 : rvCrc[4] <= 32'h736f20fa;
8'hd8 : rvCrc[4] <= 32'hc9650ce8;
8'hd9 : rvCrc[4] <= 32'h80686b65;
8'hda : rvCrc[4] <= 32'h5b7fc3f2;
8'hdb : rvCrc[4] <= 32'h1272a47f;
8'hdc : rvCrc[4] <= 32'he9918f6b;
8'hdd : rvCrc[4] <= 32'ha09ce8e6;
8'hde : rvCrc[4] <= 32'h7b8b4071;
8'hdf : rvCrc[4] <= 32'h328627fc;
8'he0 : rvCrc[4] <= 32'h083b044d;
8'he1 : rvCrc[4] <= 32'h413663c0;
8'he2 : rvCrc[4] <= 32'h9a21cb57;
8'he3 : rvCrc[4] <= 32'hd32cacda;
8'he4 : rvCrc[4] <= 32'h28cf87ce;
8'he5 : rvCrc[4] <= 32'h61c2e043;
8'he6 : rvCrc[4] <= 32'hbad548d4;
8'he7 : rvCrc[4] <= 32'hf3d82f59;
8'he8 : rvCrc[4] <= 32'h49d2034b;
8'he9 : rvCrc[4] <= 32'h00df64c6;
8'hea : rvCrc[4] <= 32'hdbc8cc51;
8'heb : rvCrc[4] <= 32'h92c5abdc;
8'hec : rvCrc[4] <= 32'h692680c8;
8'hed : rvCrc[4] <= 32'h202be745;
8'hee : rvCrc[4] <= 32'hfb3c4fd2;
8'hef : rvCrc[4] <= 32'hb231285f;
8'hf0 : rvCrc[4] <= 32'h8be90a41;
8'hf1 : rvCrc[4] <= 32'hc2e46dcc;
8'hf2 : rvCrc[4] <= 32'h19f3c55b;
8'hf3 : rvCrc[4] <= 32'h50fea2d6;
8'hf4 : rvCrc[4] <= 32'hab1d89c2;
8'hf5 : rvCrc[4] <= 32'he210ee4f;
8'hf6 : rvCrc[4] <= 32'h390746d8;
8'hf7 : rvCrc[4] <= 32'h700a2155;
8'hf8 : rvCrc[4] <= 32'hca000d47;
8'hf9 : rvCrc[4] <= 32'h830d6aca;
8'hfa : rvCrc[4] <= 32'h581ac25d;
8'hfb : rvCrc[4] <= 32'h1117a5d0;
8'hfc : rvCrc[4] <= 32'heaf48ec4;
8'hfd : rvCrc[4] <= 32'ha3f9e949;
8'hfe : rvCrc[4] <= 32'h78ee41de;
8'hff : rvCrc[4] <= 32'h31e32653;
endcase
case(iv_Input[047:040])
8'h00 : rvCrc[5] <= 32'h00000000;
8'h01 : rvCrc[5] <= 32'h1b280d78;
8'h02 : rvCrc[5] <= 32'h36501af0;
8'h03 : rvCrc[5] <= 32'h2d781788;
8'h04 : rvCrc[5] <= 32'h6ca035e0;
8'h05 : rvCrc[5] <= 32'h77883898;
8'h06 : rvCrc[5] <= 32'h5af02f10;
8'h07 : rvCrc[5] <= 32'h41d82268;
8'h08 : rvCrc[5] <= 32'hd9406bc0;
8'h09 : rvCrc[5] <= 32'hc26866b8;
8'h0a : rvCrc[5] <= 32'hef107130;
8'h0b : rvCrc[5] <= 32'hf4387c48;
8'h0c : rvCrc[5] <= 32'hb5e05e20;
8'h0d : rvCrc[5] <= 32'haec85358;
8'h0e : rvCrc[5] <= 32'h83b044d0;
8'h0f : rvCrc[5] <= 32'h989849a8;
8'h10 : rvCrc[5] <= 32'hb641ca37;
8'h11 : rvCrc[5] <= 32'had69c74f;
8'h12 : rvCrc[5] <= 32'h8011d0c7;
8'h13 : rvCrc[5] <= 32'h9b39ddbf;
8'h14 : rvCrc[5] <= 32'hdae1ffd7;
8'h15 : rvCrc[5] <= 32'hc1c9f2af;
8'h16 : rvCrc[5] <= 32'hecb1e527;
8'h17 : rvCrc[5] <= 32'hf799e85f;
8'h18 : rvCrc[5] <= 32'h6f01a1f7;
8'h19 : rvCrc[5] <= 32'h7429ac8f;
8'h1a : rvCrc[5] <= 32'h5951bb07;
8'h1b : rvCrc[5] <= 32'h4279b67f;
8'h1c : rvCrc[5] <= 32'h03a19417;
8'h1d : rvCrc[5] <= 32'h1889996f;
8'h1e : rvCrc[5] <= 32'h35f18ee7;
8'h1f : rvCrc[5] <= 32'h2ed9839f;
8'h20 : rvCrc[5] <= 32'h684289d9;
8'h21 : rvCrc[5] <= 32'h736a84a1;
8'h22 : rvCrc[5] <= 32'h5e129329;
8'h23 : rvCrc[5] <= 32'h453a9e51;
8'h24 : rvCrc[5] <= 32'h04e2bc39;
8'h25 : rvCrc[5] <= 32'h1fcab141;
8'h26 : rvCrc[5] <= 32'h32b2a6c9;
8'h27 : rvCrc[5] <= 32'h299aabb1;
8'h28 : rvCrc[5] <= 32'hb102e219;
8'h29 : rvCrc[5] <= 32'haa2aef61;
8'h2a : rvCrc[5] <= 32'h8752f8e9;
8'h2b : rvCrc[5] <= 32'h9c7af591;
8'h2c : rvCrc[5] <= 32'hdda2d7f9;
8'h2d : rvCrc[5] <= 32'hc68ada81;
8'h2e : rvCrc[5] <= 32'hebf2cd09;
8'h2f : rvCrc[5] <= 32'hf0dac071;
8'h30 : rvCrc[5] <= 32'hde0343ee;
8'h31 : rvCrc[5] <= 32'hc52b4e96;
8'h32 : rvCrc[5] <= 32'he853591e;
8'h33 : rvCrc[5] <= 32'hf37b5466;
8'h34 : rvCrc[5] <= 32'hb2a3760e;
8'h35 : rvCrc[5] <= 32'ha98b7b76;
8'h36 : rvCrc[5] <= 32'h84f36cfe;
8'h37 : rvCrc[5] <= 32'h9fdb6186;
8'h38 : rvCrc[5] <= 32'h0743282e;
8'h39 : rvCrc[5] <= 32'h1c6b2556;
8'h3a : rvCrc[5] <= 32'h311332de;
8'h3b : rvCrc[5] <= 32'h2a3b3fa6;
8'h3c : rvCrc[5] <= 32'h6be31dce;
8'h3d : rvCrc[5] <= 32'h70cb10b6;
8'h3e : rvCrc[5] <= 32'h5db3073e;
8'h3f : rvCrc[5] <= 32'h469b0a46;
8'h40 : rvCrc[5] <= 32'hd08513b2;
8'h41 : rvCrc[5] <= 32'hcbad1eca;
8'h42 : rvCrc[5] <= 32'he6d50942;
8'h43 : rvCrc[5] <= 32'hfdfd043a;
8'h44 : rvCrc[5] <= 32'hbc252652;
8'h45 : rvCrc[5] <= 32'ha70d2b2a;
8'h46 : rvCrc[5] <= 32'h8a753ca2;
8'h47 : rvCrc[5] <= 32'h915d31da;
8'h48 : rvCrc[5] <= 32'h09c57872;
8'h49 : rvCrc[5] <= 32'h12ed750a;
8'h4a : rvCrc[5] <= 32'h3f956282;
8'h4b : rvCrc[5] <= 32'h24bd6ffa;
8'h4c : rvCrc[5] <= 32'h65654d92;
8'h4d : rvCrc[5] <= 32'h7e4d40ea;
8'h4e : rvCrc[5] <= 32'h53355762;
8'h4f : rvCrc[5] <= 32'h481d5a1a;
8'h50 : rvCrc[5] <= 32'h66c4d985;
8'h51 : rvCrc[5] <= 32'h7decd4fd;
8'h52 : rvCrc[5] <= 32'h5094c375;
8'h53 : rvCrc[5] <= 32'h4bbcce0d;
8'h54 : rvCrc[5] <= 32'h0a64ec65;
8'h55 : rvCrc[5] <= 32'h114ce11d;
8'h56 : rvCrc[5] <= 32'h3c34f695;
8'h57 : rvCrc[5] <= 32'h271cfbed;
8'h58 : rvCrc[5] <= 32'hbf84b245;
8'h59 : rvCrc[5] <= 32'ha4acbf3d;
8'h5a : rvCrc[5] <= 32'h89d4a8b5;
8'h5b : rvCrc[5] <= 32'h92fca5cd;
8'h5c : rvCrc[5] <= 32'hd32487a5;
8'h5d : rvCrc[5] <= 32'hc80c8add;
8'h5e : rvCrc[5] <= 32'he5749d55;
8'h5f : rvCrc[5] <= 32'hfe5c902d;
8'h60 : rvCrc[5] <= 32'hb8c79a6b;
8'h61 : rvCrc[5] <= 32'ha3ef9713;
8'h62 : rvCrc[5] <= 32'h8e97809b;
8'h63 : rvCrc[5] <= 32'h95bf8de3;
8'h64 : rvCrc[5] <= 32'hd467af8b;
8'h65 : rvCrc[5] <= 32'hcf4fa2f3;
8'h66 : rvCrc[5] <= 32'he237b57b;
8'h67 : rvCrc[5] <= 32'hf91fb803;
8'h68 : rvCrc[5] <= 32'h6187f1ab;
8'h69 : rvCrc[5] <= 32'h7aaffcd3;
8'h6a : rvCrc[5] <= 32'h57d7eb5b;
8'h6b : rvCrc[5] <= 32'h4cffe623;
8'h6c : rvCrc[5] <= 32'h0d27c44b;
8'h6d : rvCrc[5] <= 32'h160fc933;
8'h6e : rvCrc[5] <= 32'h3b77debb;
8'h6f : rvCrc[5] <= 32'h205fd3c3;
8'h70 : rvCrc[5] <= 32'h0e86505c;
8'h71 : rvCrc[5] <= 32'h15ae5d24;
8'h72 : rvCrc[5] <= 32'h38d64aac;
8'h73 : rvCrc[5] <= 32'h23fe47d4;
8'h74 : rvCrc[5] <= 32'h622665bc;
8'h75 : rvCrc[5] <= 32'h790e68c4;
8'h76 : rvCrc[5] <= 32'h54767f4c;
8'h77 : rvCrc[5] <= 32'h4f5e7234;
8'h78 : rvCrc[5] <= 32'hd7c63b9c;
8'h79 : rvCrc[5] <= 32'hccee36e4;
8'h7a : rvCrc[5] <= 32'he196216c;
8'h7b : rvCrc[5] <= 32'hfabe2c14;
8'h7c : rvCrc[5] <= 32'hbb660e7c;
8'h7d : rvCrc[5] <= 32'ha04e0304;
8'h7e : rvCrc[5] <= 32'h8d36148c;
8'h7f : rvCrc[5] <= 32'h961e19f4;
8'h80 : rvCrc[5] <= 32'ha5cb3ad3;
8'h81 : rvCrc[5] <= 32'hbee337ab;
8'h82 : rvCrc[5] <= 32'h939b2023;
8'h83 : rvCrc[5] <= 32'h88b32d5b;
8'h84 : rvCrc[5] <= 32'hc96b0f33;
8'h85 : rvCrc[5] <= 32'hd243024b;
8'h86 : rvCrc[5] <= 32'hff3b15c3;
8'h87 : rvCrc[5] <= 32'he41318bb;
8'h88 : rvCrc[5] <= 32'h7c8b5113;
8'h89 : rvCrc[5] <= 32'h67a35c6b;
8'h8a : rvCrc[5] <= 32'h4adb4be3;
8'h8b : rvCrc[5] <= 32'h51f3469b;
8'h8c : rvCrc[5] <= 32'h102b64f3;
8'h8d : rvCrc[5] <= 32'h0b03698b;
8'h8e : rvCrc[5] <= 32'h267b7e03;
8'h8f : rvCrc[5] <= 32'h3d53737b;
8'h90 : rvCrc[5] <= 32'h138af0e4;
8'h91 : rvCrc[5] <= 32'h08a2fd9c;
8'h92 : rvCrc[5] <= 32'h25daea14;
8'h93 : rvCrc[5] <= 32'h3ef2e76c;
8'h94 : rvCrc[5] <= 32'h7f2ac504;
8'h95 : rvCrc[5] <= 32'h6402c87c;
8'h96 : rvCrc[5] <= 32'h497adff4;
8'h97 : rvCrc[5] <= 32'h5252d28c;
8'h98 : rvCrc[5] <= 32'hcaca9b24;
8'h99 : rvCrc[5] <= 32'hd1e2965c;
8'h9a : rvCrc[5] <= 32'hfc9a81d4;
8'h9b : rvCrc[5] <= 32'he7b28cac;
8'h9c : rvCrc[5] <= 32'ha66aaec4;
8'h9d : rvCrc[5] <= 32'hbd42a3bc;
8'h9e : rvCrc[5] <= 32'h903ab434;
8'h9f : rvCrc[5] <= 32'h8b12b94c;
8'ha0 : rvCrc[5] <= 32'hcd89b30a;
8'ha1 : rvCrc[5] <= 32'hd6a1be72;
8'ha2 : rvCrc[5] <= 32'hfbd9a9fa;
8'ha3 : rvCrc[5] <= 32'he0f1a482;
8'ha4 : rvCrc[5] <= 32'ha12986ea;
8'ha5 : rvCrc[5] <= 32'hba018b92;
8'ha6 : rvCrc[5] <= 32'h97799c1a;
8'ha7 : rvCrc[5] <= 32'h8c519162;
8'ha8 : rvCrc[5] <= 32'h14c9d8ca;
8'ha9 : rvCrc[5] <= 32'h0fe1d5b2;
8'haa : rvCrc[5] <= 32'h2299c23a;
8'hab : rvCrc[5] <= 32'h39b1cf42;
8'hac : rvCrc[5] <= 32'h7869ed2a;
8'had : rvCrc[5] <= 32'h6341e052;
8'hae : rvCrc[5] <= 32'h4e39f7da;
8'haf : rvCrc[5] <= 32'h5511faa2;
8'hb0 : rvCrc[5] <= 32'h7bc8793d;
8'hb1 : rvCrc[5] <= 32'h60e07445;
8'hb2 : rvCrc[5] <= 32'h4d9863cd;
8'hb3 : rvCrc[5] <= 32'h56b06eb5;
8'hb4 : rvCrc[5] <= 32'h17684cdd;
8'hb5 : rvCrc[5] <= 32'h0c4041a5;
8'hb6 : rvCrc[5] <= 32'h2138562d;
8'hb7 : rvCrc[5] <= 32'h3a105b55;
8'hb8 : rvCrc[5] <= 32'ha28812fd;
8'hb9 : rvCrc[5] <= 32'hb9a01f85;
8'hba : rvCrc[5] <= 32'h94d8080d;
8'hbb : rvCrc[5] <= 32'h8ff00575;
8'hbc : rvCrc[5] <= 32'hce28271d;
8'hbd : rvCrc[5] <= 32'hd5002a65;
8'hbe : rvCrc[5] <= 32'hf8783ded;
8'hbf : rvCrc[5] <= 32'he3503095;
8'hc0 : rvCrc[5] <= 32'h754e2961;
8'hc1 : rvCrc[5] <= 32'h6e662419;
8'hc2 : rvCrc[5] <= 32'h431e3391;
8'hc3 : rvCrc[5] <= 32'h58363ee9;
8'hc4 : rvCrc[5] <= 32'h19ee1c81;
8'hc5 : rvCrc[5] <= 32'h02c611f9;
8'hc6 : rvCrc[5] <= 32'h2fbe0671;
8'hc7 : rvCrc[5] <= 32'h34960b09;
8'hc8 : rvCrc[5] <= 32'hac0e42a1;
8'hc9 : rvCrc[5] <= 32'hb7264fd9;
8'hca : rvCrc[5] <= 32'h9a5e5851;
8'hcb : rvCrc[5] <= 32'h81765529;
8'hcc : rvCrc[5] <= 32'hc0ae7741;
8'hcd : rvCrc[5] <= 32'hdb867a39;
8'hce : rvCrc[5] <= 32'hf6fe6db1;
8'hcf : rvCrc[5] <= 32'hedd660c9;
8'hd0 : rvCrc[5] <= 32'hc30fe356;
8'hd1 : rvCrc[5] <= 32'hd827ee2e;
8'hd2 : rvCrc[5] <= 32'hf55ff9a6;
8'hd3 : rvCrc[5] <= 32'hee77f4de;
8'hd4 : rvCrc[5] <= 32'hafafd6b6;
8'hd5 : rvCrc[5] <= 32'hb487dbce;
8'hd6 : rvCrc[5] <= 32'h99ffcc46;
8'hd7 : rvCrc[5] <= 32'h82d7c13e;
8'hd8 : rvCrc[5] <= 32'h1a4f8896;
8'hd9 : rvCrc[5] <= 32'h016785ee;
8'hda : rvCrc[5] <= 32'h2c1f9266;
8'hdb : rvCrc[5] <= 32'h37379f1e;
8'hdc : rvCrc[5] <= 32'h76efbd76;
8'hdd : rvCrc[5] <= 32'h6dc7b00e;
8'hde : rvCrc[5] <= 32'h40bfa786;
8'hdf : rvCrc[5] <= 32'h5b97aafe;
8'he0 : rvCrc[5] <= 32'h1d0ca0b8;
8'he1 : rvCrc[5] <= 32'h0624adc0;
8'he2 : rvCrc[5] <= 32'h2b5cba48;
8'he3 : rvCrc[5] <= 32'h3074b730;
8'he4 : rvCrc[5] <= 32'h71ac9558;
8'he5 : rvCrc[5] <= 32'h6a849820;
8'he6 : rvCrc[5] <= 32'h47fc8fa8;
8'he7 : rvCrc[5] <= 32'h5cd482d0;
8'he8 : rvCrc[5] <= 32'hc44ccb78;
8'he9 : rvCrc[5] <= 32'hdf64c600;
8'hea : rvCrc[5] <= 32'hf21cd188;
8'heb : rvCrc[5] <= 32'he934dcf0;
8'hec : rvCrc[5] <= 32'ha8ecfe98;
8'hed : rvCrc[5] <= 32'hb3c4f3e0;
8'hee : rvCrc[5] <= 32'h9ebce468;
8'hef : rvCrc[5] <= 32'h8594e910;
8'hf0 : rvCrc[5] <= 32'hab4d6a8f;
8'hf1 : rvCrc[5] <= 32'hb06567f7;
8'hf2 : rvCrc[5] <= 32'h9d1d707f;
8'hf3 : rvCrc[5] <= 32'h86357d07;
8'hf4 : rvCrc[5] <= 32'hc7ed5f6f;
8'hf5 : rvCrc[5] <= 32'hdcc55217;
8'hf6 : rvCrc[5] <= 32'hf1bd459f;
8'hf7 : rvCrc[5] <= 32'hea9548e7;
8'hf8 : rvCrc[5] <= 32'h720d014f;
8'hf9 : rvCrc[5] <= 32'h69250c37;
8'hfa : rvCrc[5] <= 32'h445d1bbf;
8'hfb : rvCrc[5] <= 32'h5f7516c7;
8'hfc : rvCrc[5] <= 32'h1ead34af;
8'hfd : rvCrc[5] <= 32'h058539d7;
8'hfe : rvCrc[5] <= 32'h28fd2e5f;
8'hff : rvCrc[5] <= 32'h33d52327;
endcase
case(iv_Input[055:048])
8'h00 : rvCrc[6] <= 32'h00000000;
8'h01 : rvCrc[6] <= 32'h4f576811;
8'h02 : rvCrc[6] <= 32'h9eaed022;
8'h03 : rvCrc[6] <= 32'hd1f9b833;
8'h04 : rvCrc[6] <= 32'h399cbdf3;
8'h05 : rvCrc[6] <= 32'h76cbd5e2;
8'h06 : rvCrc[6] <= 32'ha7326dd1;
8'h07 : rvCrc[6] <= 32'he86505c0;
8'h08 : rvCrc[6] <= 32'h73397be6;
8'h09 : rvCrc[6] <= 32'h3c6e13f7;
8'h0a : rvCrc[6] <= 32'hed97abc4;
8'h0b : rvCrc[6] <= 32'ha2c0c3d5;
8'h0c : rvCrc[6] <= 32'h4aa5c615;
8'h0d : rvCrc[6] <= 32'h05f2ae04;
8'h0e : rvCrc[6] <= 32'hd40b1637;
8'h0f : rvCrc[6] <= 32'h9b5c7e26;
8'h10 : rvCrc[6] <= 32'he672f7cc;
8'h11 : rvCrc[6] <= 32'ha9259fdd;
8'h12 : rvCrc[6] <= 32'h78dc27ee;
8'h13 : rvCrc[6] <= 32'h378b4fff;
8'h14 : rvCrc[6] <= 32'hdfee4a3f;
8'h15 : rvCrc[6] <= 32'h90b9222e;
8'h16 : rvCrc[6] <= 32'h41409a1d;
8'h17 : rvCrc[6] <= 32'h0e17f20c;
8'h18 : rvCrc[6] <= 32'h954b8c2a;
8'h19 : rvCrc[6] <= 32'hda1ce43b;
8'h1a : rvCrc[6] <= 32'h0be55c08;
8'h1b : rvCrc[6] <= 32'h44b23419;
8'h1c : rvCrc[6] <= 32'hacd731d9;
8'h1d : rvCrc[6] <= 32'he38059c8;
8'h1e : rvCrc[6] <= 32'h3279e1fb;
8'h1f : rvCrc[6] <= 32'h7d2e89ea;
8'h20 : rvCrc[6] <= 32'hc824f22f;
8'h21 : rvCrc[6] <= 32'h87739a3e;
8'h22 : rvCrc[6] <= 32'h568a220d;
8'h23 : rvCrc[6] <= 32'h19dd4a1c;
8'h24 : rvCrc[6] <= 32'hf1b84fdc;
8'h25 : rvCrc[6] <= 32'hbeef27cd;
8'h26 : rvCrc[6] <= 32'h6f169ffe;
8'h27 : rvCrc[6] <= 32'h2041f7ef;
8'h28 : rvCrc[6] <= 32'hbb1d89c9;
8'h29 : rvCrc[6] <= 32'hf44ae1d8;
8'h2a : rvCrc[6] <= 32'h25b359eb;
8'h2b : rvCrc[6] <= 32'h6ae431fa;
8'h2c : rvCrc[6] <= 32'h8281343a;
8'h2d : rvCrc[6] <= 32'hcdd65c2b;
8'h2e : rvCrc[6] <= 32'h1c2fe418;
8'h2f : rvCrc[6] <= 32'h53788c09;
8'h30 : rvCrc[6] <= 32'h2e5605e3;
8'h31 : rvCrc[6] <= 32'h61016df2;
8'h32 : rvCrc[6] <= 32'hb0f8d5c1;
8'h33 : rvCrc[6] <= 32'hffafbdd0;
8'h34 : rvCrc[6] <= 32'h17cab810;
8'h35 : rvCrc[6] <= 32'h589dd001;
8'h36 : rvCrc[6] <= 32'h89646832;
8'h37 : rvCrc[6] <= 32'hc6330023;
8'h38 : rvCrc[6] <= 32'h5d6f7e05;
8'h39 : rvCrc[6] <= 32'h12381614;
8'h3a : rvCrc[6] <= 32'hc3c1ae27;
8'h3b : rvCrc[6] <= 32'h8c96c636;
8'h3c : rvCrc[6] <= 32'h64f3c3f6;
8'h3d : rvCrc[6] <= 32'h2ba4abe7;
8'h3e : rvCrc[6] <= 32'hfa5d13d4;
8'h3f : rvCrc[6] <= 32'hb50a7bc5;
8'h40 : rvCrc[6] <= 32'h9488f9e9;
8'h41 : rvCrc[6] <= 32'hdbdf91f8;
8'h42 : rvCrc[6] <= 32'h0a2629cb;
8'h43 : rvCrc[6] <= 32'h457141da;
8'h44 : rvCrc[6] <= 32'had14441a;
8'h45 : rvCrc[6] <= 32'he2432c0b;
8'h46 : rvCrc[6] <= 32'h33ba9438;
8'h47 : rvCrc[6] <= 32'h7cedfc29;
8'h48 : rvCrc[6] <= 32'he7b1820f;
8'h49 : rvCrc[6] <= 32'ha8e6ea1e;
8'h4a : rvCrc[6] <= 32'h791f522d;
8'h4b : rvCrc[6] <= 32'h36483a3c;
8'h4c : rvCrc[6] <= 32'hde2d3ffc;
8'h4d : rvCrc[6] <= 32'h917a57ed;
8'h4e : rvCrc[6] <= 32'h4083efde;
8'h4f : rvCrc[6] <= 32'h0fd487cf;
8'h50 : rvCrc[6] <= 32'h72fa0e25;
8'h51 : rvCrc[6] <= 32'h3dad6634;
8'h52 : rvCrc[6] <= 32'hec54de07;
8'h53 : rvCrc[6] <= 32'ha303b616;
8'h54 : rvCrc[6] <= 32'h4b66b3d6;
8'h55 : rvCrc[6] <= 32'h0431dbc7;
8'h56 : rvCrc[6] <= 32'hd5c863f4;
8'h57 : rvCrc[6] <= 32'h9a9f0be5;
8'h58 : rvCrc[6] <= 32'h01c375c3;
8'h59 : rvCrc[6] <= 32'h4e941dd2;
8'h5a : rvCrc[6] <= 32'h9f6da5e1;
8'h5b : rvCrc[6] <= 32'hd03acdf0;
8'h5c : rvCrc[6] <= 32'h385fc830;
8'h5d : rvCrc[6] <= 32'h7708a021;
8'h5e : rvCrc[6] <= 32'ha6f11812;
8'h5f : rvCrc[6] <= 32'he9a67003;
8'h60 : rvCrc[6] <= 32'h5cac0bc6;
8'h61 : rvCrc[6] <= 32'h13fb63d7;
8'h62 : rvCrc[6] <= 32'hc202dbe4;
8'h63 : rvCrc[6] <= 32'h8d55b3f5;
8'h64 : rvCrc[6] <= 32'h6530b635;
8'h65 : rvCrc[6] <= 32'h2a67de24;
8'h66 : rvCrc[6] <= 32'hfb9e6617;
8'h67 : rvCrc[6] <= 32'hb4c90e06;
8'h68 : rvCrc[6] <= 32'h2f957020;
8'h69 : rvCrc[6] <= 32'h60c21831;
8'h6a : rvCrc[6] <= 32'hb13ba002;
8'h6b : rvCrc[6] <= 32'hfe6cc813;
8'h6c : rvCrc[6] <= 32'h1609cdd3;
8'h6d : rvCrc[6] <= 32'h595ea5c2;
8'h6e : rvCrc[6] <= 32'h88a71df1;
8'h6f : rvCrc[6] <= 32'hc7f075e0;
8'h70 : rvCrc[6] <= 32'hbadefc0a;
8'h71 : rvCrc[6] <= 32'hf589941b;
8'h72 : rvCrc[6] <= 32'h24702c28;
8'h73 : rvCrc[6] <= 32'h6b274439;
8'h74 : rvCrc[6] <= 32'h834241f9;
8'h75 : rvCrc[6] <= 32'hcc1529e8;
8'h76 : rvCrc[6] <= 32'h1dec91db;
8'h77 : rvCrc[6] <= 32'h52bbf9ca;
8'h78 : rvCrc[6] <= 32'hc9e787ec;
8'h79 : rvCrc[6] <= 32'h86b0effd;
8'h7a : rvCrc[6] <= 32'h574957ce;
8'h7b : rvCrc[6] <= 32'h181e3fdf;
8'h7c : rvCrc[6] <= 32'hf07b3a1f;
8'h7d : rvCrc[6] <= 32'hbf2c520e;
8'h7e : rvCrc[6] <= 32'h6ed5ea3d;
8'h7f : rvCrc[6] <= 32'h2182822c;
8'h80 : rvCrc[6] <= 32'h2dd0ee65;
8'h81 : rvCrc[6] <= 32'h62878674;
8'h82 : rvCrc[6] <= 32'hb37e3e47;
8'h83 : rvCrc[6] <= 32'hfc295656;
8'h84 : rvCrc[6] <= 32'h144c5396;
8'h85 : rvCrc[6] <= 32'h5b1b3b87;
8'h86 : rvCrc[6] <= 32'h8ae283b4;
8'h87 : rvCrc[6] <= 32'hc5b5eba5;
8'h88 : rvCrc[6] <= 32'h5ee99583;
8'h89 : rvCrc[6] <= 32'h11befd92;
8'h8a : rvCrc[6] <= 32'hc04745a1;
8'h8b : rvCrc[6] <= 32'h8f102db0;
8'h8c : rvCrc[6] <= 32'h67752870;
8'h8d : rvCrc[6] <= 32'h28224061;
8'h8e : rvCrc[6] <= 32'hf9dbf852;
8'h8f : rvCrc[6] <= 32'hb68c9043;
8'h90 : rvCrc[6] <= 32'hcba219a9;
8'h91 : rvCrc[6] <= 32'h84f571b8;
8'h92 : rvCrc[6] <= 32'h550cc98b;
8'h93 : rvCrc[6] <= 32'h1a5ba19a;
8'h94 : rvCrc[6] <= 32'hf23ea45a;
8'h95 : rvCrc[6] <= 32'hbd69cc4b;
8'h96 : rvCrc[6] <= 32'h6c907478;
8'h97 : rvCrc[6] <= 32'h23c71c69;
8'h98 : rvCrc[6] <= 32'hb89b624f;
8'h99 : rvCrc[6] <= 32'hf7cc0a5e;
8'h9a : rvCrc[6] <= 32'h2635b26d;
8'h9b : rvCrc[6] <= 32'h6962da7c;
8'h9c : rvCrc[6] <= 32'h8107dfbc;
8'h9d : rvCrc[6] <= 32'hce50b7ad;
8'h9e : rvCrc[6] <= 32'h1fa90f9e;
8'h9f : rvCrc[6] <= 32'h50fe678f;
8'ha0 : rvCrc[6] <= 32'he5f41c4a;
8'ha1 : rvCrc[6] <= 32'haaa3745b;
8'ha2 : rvCrc[6] <= 32'h7b5acc68;
8'ha3 : rvCrc[6] <= 32'h340da479;
8'ha4 : rvCrc[6] <= 32'hdc68a1b9;
8'ha5 : rvCrc[6] <= 32'h933fc9a8;
8'ha6 : rvCrc[6] <= 32'h42c6719b;
8'ha7 : rvCrc[6] <= 32'h0d91198a;
8'ha8 : rvCrc[6] <= 32'h96cd67ac;
8'ha9 : rvCrc[6] <= 32'hd99a0fbd;
8'haa : rvCrc[6] <= 32'h0863b78e;
8'hab : rvCrc[6] <= 32'h4734df9f;
8'hac : rvCrc[6] <= 32'haf51da5f;
8'had : rvCrc[6] <= 32'he006b24e;
8'hae : rvCrc[6] <= 32'h31ff0a7d;
8'haf : rvCrc[6] <= 32'h7ea8626c;
8'hb0 : rvCrc[6] <= 32'h0386eb86;
8'hb1 : rvCrc[6] <= 32'h4cd18397;
8'hb2 : rvCrc[6] <= 32'h9d283ba4;
8'hb3 : rvCrc[6] <= 32'hd27f53b5;
8'hb4 : rvCrc[6] <= 32'h3a1a5675;
8'hb5 : rvCrc[6] <= 32'h754d3e64;
8'hb6 : rvCrc[6] <= 32'ha4b48657;
8'hb7 : rvCrc[6] <= 32'hebe3ee46;
8'hb8 : rvCrc[6] <= 32'h70bf9060;
8'hb9 : rvCrc[6] <= 32'h3fe8f871;
8'hba : rvCrc[6] <= 32'hee114042;
8'hbb : rvCrc[6] <= 32'ha1462853;
8'hbc : rvCrc[6] <= 32'h49232d93;
8'hbd : rvCrc[6] <= 32'h06744582;
8'hbe : rvCrc[6] <= 32'hd78dfdb1;
8'hbf : rvCrc[6] <= 32'h98da95a0;
8'hc0 : rvCrc[6] <= 32'hb958178c;
8'hc1 : rvCrc[6] <= 32'hf60f7f9d;
8'hc2 : rvCrc[6] <= 32'h27f6c7ae;
8'hc3 : rvCrc[6] <= 32'h68a1afbf;
8'hc4 : rvCrc[6] <= 32'h80c4aa7f;
8'hc5 : rvCrc[6] <= 32'hcf93c26e;
8'hc6 : rvCrc[6] <= 32'h1e6a7a5d;
8'hc7 : rvCrc[6] <= 32'h513d124c;
8'hc8 : rvCrc[6] <= 32'hca616c6a;
8'hc9 : rvCrc[6] <= 32'h8536047b;
8'hca : rvCrc[6] <= 32'h54cfbc48;
8'hcb : rvCrc[6] <= 32'h1b98d459;
8'hcc : rvCrc[6] <= 32'hf3fdd199;
8'hcd : rvCrc[6] <= 32'hbcaab988;
8'hce : rvCrc[6] <= 32'h6d5301bb;
8'hcf : rvCrc[6] <= 32'h220469aa;
8'hd0 : rvCrc[6] <= 32'h5f2ae040;
8'hd1 : rvCrc[6] <= 32'h107d8851;
8'hd2 : rvCrc[6] <= 32'hc1843062;
8'hd3 : rvCrc[6] <= 32'h8ed35873;
8'hd4 : rvCrc[6] <= 32'h66b65db3;
8'hd5 : rvCrc[6] <= 32'h29e135a2;
8'hd6 : rvCrc[6] <= 32'hf8188d91;
8'hd7 : rvCrc[6] <= 32'hb74fe580;
8'hd8 : rvCrc[6] <= 32'h2c139ba6;
8'hd9 : rvCrc[6] <= 32'h6344f3b7;
8'hda : rvCrc[6] <= 32'hb2bd4b84;
8'hdb : rvCrc[6] <= 32'hfdea2395;
8'hdc : rvCrc[6] <= 32'h158f2655;
8'hdd : rvCrc[6] <= 32'h5ad84e44;
8'hde : rvCrc[6] <= 32'h8b21f677;
8'hdf : rvCrc[6] <= 32'hc4769e66;
8'he0 : rvCrc[6] <= 32'h717ce5a3;
8'he1 : rvCrc[6] <= 32'h3e2b8db2;
8'he2 : rvCrc[6] <= 32'hefd23581;
8'he3 : rvCrc[6] <= 32'ha0855d90;
8'he4 : rvCrc[6] <= 32'h48e05850;
8'he5 : rvCrc[6] <= 32'h07b73041;
8'he6 : rvCrc[6] <= 32'hd64e8872;
8'he7 : rvCrc[6] <= 32'h9919e063;
8'he8 : rvCrc[6] <= 32'h02459e45;
8'he9 : rvCrc[6] <= 32'h4d12f654;
8'hea : rvCrc[6] <= 32'h9ceb4e67;
8'heb : rvCrc[6] <= 32'hd3bc2676;
8'hec : rvCrc[6] <= 32'h3bd923b6;
8'hed : rvCrc[6] <= 32'h748e4ba7;
8'hee : rvCrc[6] <= 32'ha577f394;
8'hef : rvCrc[6] <= 32'hea209b85;
8'hf0 : rvCrc[6] <= 32'h970e126f;
8'hf1 : rvCrc[6] <= 32'hd8597a7e;
8'hf2 : rvCrc[6] <= 32'h09a0c24d;
8'hf3 : rvCrc[6] <= 32'h46f7aa5c;
8'hf4 : rvCrc[6] <= 32'hae92af9c;
8'hf5 : rvCrc[6] <= 32'he1c5c78d;
8'hf6 : rvCrc[6] <= 32'h303c7fbe;
8'hf7 : rvCrc[6] <= 32'h7f6b17af;
8'hf8 : rvCrc[6] <= 32'he4376989;
8'hf9 : rvCrc[6] <= 32'hab600198;
8'hfa : rvCrc[6] <= 32'h7a99b9ab;
8'hfb : rvCrc[6] <= 32'h35ced1ba;
8'hfc : rvCrc[6] <= 32'hddabd47a;
8'hfd : rvCrc[6] <= 32'h92fcbc6b;
8'hfe : rvCrc[6] <= 32'h43050458;
8'hff : rvCrc[6] <= 32'h0c526c49;
endcase
case(iv_Input[063:056])
8'h00 : rvCrc[7] <= 32'h00000000;
8'h01 : rvCrc[7] <= 32'h5ba1dcca;
8'h02 : rvCrc[7] <= 32'hb743b994;
8'h03 : rvCrc[7] <= 32'hece2655e;
8'h04 : rvCrc[7] <= 32'h6a466e9f;
8'h05 : rvCrc[7] <= 32'h31e7b255;
8'h06 : rvCrc[7] <= 32'hdd05d70b;
8'h07 : rvCrc[7] <= 32'h86a40bc1;
8'h08 : rvCrc[7] <= 32'hd48cdd3e;
8'h09 : rvCrc[7] <= 32'h8f2d01f4;
8'h0a : rvCrc[7] <= 32'h63cf64aa;
8'h0b : rvCrc[7] <= 32'h386eb860;
8'h0c : rvCrc[7] <= 32'hbecab3a1;
8'h0d : rvCrc[7] <= 32'he56b6f6b;
8'h0e : rvCrc[7] <= 32'h09890a35;
8'h0f : rvCrc[7] <= 32'h5228d6ff;
8'h10 : rvCrc[7] <= 32'hadd8a7cb;
8'h11 : rvCrc[7] <= 32'hf6797b01;
8'h12 : rvCrc[7] <= 32'h1a9b1e5f;
8'h13 : rvCrc[7] <= 32'h413ac295;
8'h14 : rvCrc[7] <= 32'hc79ec954;
8'h15 : rvCrc[7] <= 32'h9c3f159e;
8'h16 : rvCrc[7] <= 32'h70dd70c0;
8'h17 : rvCrc[7] <= 32'h2b7cac0a;
8'h18 : rvCrc[7] <= 32'h79547af5;
8'h19 : rvCrc[7] <= 32'h22f5a63f;
8'h1a : rvCrc[7] <= 32'hce17c361;
8'h1b : rvCrc[7] <= 32'h95b61fab;
8'h1c : rvCrc[7] <= 32'h1312146a;
8'h1d : rvCrc[7] <= 32'h48b3c8a0;
8'h1e : rvCrc[7] <= 32'ha451adfe;
8'h1f : rvCrc[7] <= 32'hfff07134;
8'h20 : rvCrc[7] <= 32'h5f705221;
8'h21 : rvCrc[7] <= 32'h04d18eeb;
8'h22 : rvCrc[7] <= 32'he833ebb5;
8'h23 : rvCrc[7] <= 32'hb392377f;
8'h24 : rvCrc[7] <= 32'h35363cbe;
8'h25 : rvCrc[7] <= 32'h6e97e074;
8'h26 : rvCrc[7] <= 32'h8275852a;
8'h27 : rvCrc[7] <= 32'hd9d459e0;
8'h28 : rvCrc[7] <= 32'h8bfc8f1f;
8'h29 : rvCrc[7] <= 32'hd05d53d5;
8'h2a : rvCrc[7] <= 32'h3cbf368b;
8'h2b : rvCrc[7] <= 32'h671eea41;
8'h2c : rvCrc[7] <= 32'he1bae180;
8'h2d : rvCrc[7] <= 32'hba1b3d4a;
8'h2e : rvCrc[7] <= 32'h56f95814;
8'h2f : rvCrc[7] <= 32'h0d5884de;
8'h30 : rvCrc[7] <= 32'hf2a8f5ea;
8'h31 : rvCrc[7] <= 32'ha9092920;
8'h32 : rvCrc[7] <= 32'h45eb4c7e;
8'h33 : rvCrc[7] <= 32'h1e4a90b4;
8'h34 : rvCrc[7] <= 32'h98ee9b75;
8'h35 : rvCrc[7] <= 32'hc34f47bf;
8'h36 : rvCrc[7] <= 32'h2fad22e1;
8'h37 : rvCrc[7] <= 32'h740cfe2b;
8'h38 : rvCrc[7] <= 32'h262428d4;
8'h39 : rvCrc[7] <= 32'h7d85f41e;
8'h3a : rvCrc[7] <= 32'h91679140;
8'h3b : rvCrc[7] <= 32'hcac64d8a;
8'h3c : rvCrc[7] <= 32'h4c62464b;
8'h3d : rvCrc[7] <= 32'h17c39a81;
8'h3e : rvCrc[7] <= 32'hfb21ffdf;
8'h3f : rvCrc[7] <= 32'ha0802315;
8'h40 : rvCrc[7] <= 32'hbee0a442;
8'h41 : rvCrc[7] <= 32'he5417888;
8'h42 : rvCrc[7] <= 32'h09a31dd6;
8'h43 : rvCrc[7] <= 32'h5202c11c;
8'h44 : rvCrc[7] <= 32'hd4a6cadd;
8'h45 : rvCrc[7] <= 32'h8f071617;
8'h46 : rvCrc[7] <= 32'h63e57349;
8'h47 : rvCrc[7] <= 32'h3844af83;
8'h48 : rvCrc[7] <= 32'h6a6c797c;
8'h49 : rvCrc[7] <= 32'h31cda5b6;
8'h4a : rvCrc[7] <= 32'hdd2fc0e8;
8'h4b : rvCrc[7] <= 32'h868e1c22;
8'h4c : rvCrc[7] <= 32'h002a17e3;
8'h4d : rvCrc[7] <= 32'h5b8bcb29;
8'h4e : rvCrc[7] <= 32'hb769ae77;
8'h4f : rvCrc[7] <= 32'hecc872bd;
8'h50 : rvCrc[7] <= 32'h13380389;
8'h51 : rvCrc[7] <= 32'h4899df43;
8'h52 : rvCrc[7] <= 32'ha47bba1d;
8'h53 : rvCrc[7] <= 32'hffda66d7;
8'h54 : rvCrc[7] <= 32'h797e6d16;
8'h55 : rvCrc[7] <= 32'h22dfb1dc;
8'h56 : rvCrc[7] <= 32'hce3dd482;
8'h57 : rvCrc[7] <= 32'h959c0848;
8'h58 : rvCrc[7] <= 32'hc7b4deb7;
8'h59 : rvCrc[7] <= 32'h9c15027d;
8'h5a : rvCrc[7] <= 32'h70f76723;
8'h5b : rvCrc[7] <= 32'h2b56bbe9;
8'h5c : rvCrc[7] <= 32'hadf2b028;
8'h5d : rvCrc[7] <= 32'hf6536ce2;
8'h5e : rvCrc[7] <= 32'h1ab109bc;
8'h5f : rvCrc[7] <= 32'h4110d576;
8'h60 : rvCrc[7] <= 32'he190f663;
8'h61 : rvCrc[7] <= 32'hba312aa9;
8'h62 : rvCrc[7] <= 32'h56d34ff7;
8'h63 : rvCrc[7] <= 32'h0d72933d;
8'h64 : rvCrc[7] <= 32'h8bd698fc;
8'h65 : rvCrc[7] <= 32'hd0774436;
8'h66 : rvCrc[7] <= 32'h3c952168;
8'h67 : rvCrc[7] <= 32'h6734fda2;
8'h68 : rvCrc[7] <= 32'h351c2b5d;
8'h69 : rvCrc[7] <= 32'h6ebdf797;
8'h6a : rvCrc[7] <= 32'h825f92c9;
8'h6b : rvCrc[7] <= 32'hd9fe4e03;
8'h6c : rvCrc[7] <= 32'h5f5a45c2;
8'h6d : rvCrc[7] <= 32'h04fb9908;
8'h6e : rvCrc[7] <= 32'he819fc56;
8'h6f : rvCrc[7] <= 32'hb3b8209c;
8'h70 : rvCrc[7] <= 32'h4c4851a8;
8'h71 : rvCrc[7] <= 32'h17e98d62;
8'h72 : rvCrc[7] <= 32'hfb0be83c;
8'h73 : rvCrc[7] <= 32'ha0aa34f6;
8'h74 : rvCrc[7] <= 32'h260e3f37;
8'h75 : rvCrc[7] <= 32'h7dafe3fd;
8'h76 : rvCrc[7] <= 32'h914d86a3;
8'h77 : rvCrc[7] <= 32'hcaec5a69;
8'h78 : rvCrc[7] <= 32'h98c48c96;
8'h79 : rvCrc[7] <= 32'hc365505c;
8'h7a : rvCrc[7] <= 32'h2f873502;
8'h7b : rvCrc[7] <= 32'h7426e9c8;
8'h7c : rvCrc[7] <= 32'hf282e209;
8'h7d : rvCrc[7] <= 32'ha9233ec3;
8'h7e : rvCrc[7] <= 32'h45c15b9d;
8'h7f : rvCrc[7] <= 32'h1e608757;
8'h80 : rvCrc[7] <= 32'h79005533;
8'h81 : rvCrc[7] <= 32'h22a189f9;
8'h82 : rvCrc[7] <= 32'hce43eca7;
8'h83 : rvCrc[7] <= 32'h95e2306d;
8'h84 : rvCrc[7] <= 32'h13463bac;
8'h85 : rvCrc[7] <= 32'h48e7e766;
8'h86 : rvCrc[7] <= 32'ha4058238;
8'h87 : rvCrc[7] <= 32'hffa45ef2;
8'h88 : rvCrc[7] <= 32'had8c880d;
8'h89 : rvCrc[7] <= 32'hf62d54c7;
8'h8a : rvCrc[7] <= 32'h1acf3199;
8'h8b : rvCrc[7] <= 32'h416eed53;
8'h8c : rvCrc[7] <= 32'hc7cae692;
8'h8d : rvCrc[7] <= 32'h9c6b3a58;
8'h8e : rvCrc[7] <= 32'h70895f06;
8'h8f : rvCrc[7] <= 32'h2b2883cc;
8'h90 : rvCrc[7] <= 32'hd4d8f2f8;
8'h91 : rvCrc[7] <= 32'h8f792e32;
8'h92 : rvCrc[7] <= 32'h639b4b6c;
8'h93 : rvCrc[7] <= 32'h383a97a6;
8'h94 : rvCrc[7] <= 32'hbe9e9c67;
8'h95 : rvCrc[7] <= 32'he53f40ad;
8'h96 : rvCrc[7] <= 32'h09dd25f3;
8'h97 : rvCrc[7] <= 32'h527cf939;
8'h98 : rvCrc[7] <= 32'h00542fc6;
8'h99 : rvCrc[7] <= 32'h5bf5f30c;
8'h9a : rvCrc[7] <= 32'hb7179652;
8'h9b : rvCrc[7] <= 32'hecb64a98;
8'h9c : rvCrc[7] <= 32'h6a124159;
8'h9d : rvCrc[7] <= 32'h31b39d93;
8'h9e : rvCrc[7] <= 32'hdd51f8cd;
8'h9f : rvCrc[7] <= 32'h86f02407;
8'ha0 : rvCrc[7] <= 32'h26700712;
8'ha1 : rvCrc[7] <= 32'h7dd1dbd8;
8'ha2 : rvCrc[7] <= 32'h9133be86;
8'ha3 : rvCrc[7] <= 32'hca92624c;
8'ha4 : rvCrc[7] <= 32'h4c36698d;
8'ha5 : rvCrc[7] <= 32'h1797b547;
8'ha6 : rvCrc[7] <= 32'hfb75d019;
8'ha7 : rvCrc[7] <= 32'ha0d40cd3;
8'ha8 : rvCrc[7] <= 32'hf2fcda2c;
8'ha9 : rvCrc[7] <= 32'ha95d06e6;
8'haa : rvCrc[7] <= 32'h45bf63b8;
8'hab : rvCrc[7] <= 32'h1e1ebf72;
8'hac : rvCrc[7] <= 32'h98bab4b3;
8'had : rvCrc[7] <= 32'hc31b6879;
8'hae : rvCrc[7] <= 32'h2ff90d27;
8'haf : rvCrc[7] <= 32'h7458d1ed;
8'hb0 : rvCrc[7] <= 32'h8ba8a0d9;
8'hb1 : rvCrc[7] <= 32'hd0097c13;
8'hb2 : rvCrc[7] <= 32'h3ceb194d;
8'hb3 : rvCrc[7] <= 32'h674ac587;
8'hb4 : rvCrc[7] <= 32'he1eece46;
8'hb5 : rvCrc[7] <= 32'hba4f128c;
8'hb6 : rvCrc[7] <= 32'h56ad77d2;
8'hb7 : rvCrc[7] <= 32'h0d0cab18;
8'hb8 : rvCrc[7] <= 32'h5f247de7;
8'hb9 : rvCrc[7] <= 32'h0485a12d;
8'hba : rvCrc[7] <= 32'he867c473;
8'hbb : rvCrc[7] <= 32'hb3c618b9;
8'hbc : rvCrc[7] <= 32'h35621378;
8'hbd : rvCrc[7] <= 32'h6ec3cfb2;
8'hbe : rvCrc[7] <= 32'h8221aaec;
8'hbf : rvCrc[7] <= 32'hd9807626;
8'hc0 : rvCrc[7] <= 32'hc7e0f171;
8'hc1 : rvCrc[7] <= 32'h9c412dbb;
8'hc2 : rvCrc[7] <= 32'h70a348e5;
8'hc3 : rvCrc[7] <= 32'h2b02942f;
8'hc4 : rvCrc[7] <= 32'hada69fee;
8'hc5 : rvCrc[7] <= 32'hf6074324;
8'hc6 : rvCrc[7] <= 32'h1ae5267a;
8'hc7 : rvCrc[7] <= 32'h4144fab0;
8'hc8 : rvCrc[7] <= 32'h136c2c4f;
8'hc9 : rvCrc[7] <= 32'h48cdf085;
8'hca : rvCrc[7] <= 32'ha42f95db;
8'hcb : rvCrc[7] <= 32'hff8e4911;
8'hcc : rvCrc[7] <= 32'h792a42d0;
8'hcd : rvCrc[7] <= 32'h228b9e1a;
8'hce : rvCrc[7] <= 32'hce69fb44;
8'hcf : rvCrc[7] <= 32'h95c8278e;
8'hd0 : rvCrc[7] <= 32'h6a3856ba;
8'hd1 : rvCrc[7] <= 32'h31998a70;
8'hd2 : rvCrc[7] <= 32'hdd7bef2e;
8'hd3 : rvCrc[7] <= 32'h86da33e4;
8'hd4 : rvCrc[7] <= 32'h007e3825;
8'hd5 : rvCrc[7] <= 32'h5bdfe4ef;
8'hd6 : rvCrc[7] <= 32'hb73d81b1;
8'hd7 : rvCrc[7] <= 32'hec9c5d7b;
8'hd8 : rvCrc[7] <= 32'hbeb48b84;
8'hd9 : rvCrc[7] <= 32'he515574e;
8'hda : rvCrc[7] <= 32'h09f73210;
8'hdb : rvCrc[7] <= 32'h5256eeda;
8'hdc : rvCrc[7] <= 32'hd4f2e51b;
8'hdd : rvCrc[7] <= 32'h8f5339d1;
8'hde : rvCrc[7] <= 32'h63b15c8f;
8'hdf : rvCrc[7] <= 32'h38108045;
8'he0 : rvCrc[7] <= 32'h9890a350;
8'he1 : rvCrc[7] <= 32'hc3317f9a;
8'he2 : rvCrc[7] <= 32'h2fd31ac4;
8'he3 : rvCrc[7] <= 32'h7472c60e;
8'he4 : rvCrc[7] <= 32'hf2d6cdcf;
8'he5 : rvCrc[7] <= 32'ha9771105;
8'he6 : rvCrc[7] <= 32'h4595745b;
8'he7 : rvCrc[7] <= 32'h1e34a891;
8'he8 : rvCrc[7] <= 32'h4c1c7e6e;
8'he9 : rvCrc[7] <= 32'h17bda2a4;
8'hea : rvCrc[7] <= 32'hfb5fc7fa;
8'heb : rvCrc[7] <= 32'ha0fe1b30;
8'hec : rvCrc[7] <= 32'h265a10f1;
8'hed : rvCrc[7] <= 32'h7dfbcc3b;
8'hee : rvCrc[7] <= 32'h9119a965;
8'hef : rvCrc[7] <= 32'hcab875af;
8'hf0 : rvCrc[7] <= 32'h3548049b;
8'hf1 : rvCrc[7] <= 32'h6ee9d851;
8'hf2 : rvCrc[7] <= 32'h820bbd0f;
8'hf3 : rvCrc[7] <= 32'hd9aa61c5;
8'hf4 : rvCrc[7] <= 32'h5f0e6a04;
8'hf5 : rvCrc[7] <= 32'h04afb6ce;
8'hf6 : rvCrc[7] <= 32'he84dd390;
8'hf7 : rvCrc[7] <= 32'hb3ec0f5a;
8'hf8 : rvCrc[7] <= 32'he1c4d9a5;
8'hf9 : rvCrc[7] <= 32'hba65056f;
8'hfa : rvCrc[7] <= 32'h56876031;
8'hfb : rvCrc[7] <= 32'h0d26bcfb;
8'hfc : rvCrc[7] <= 32'h8b82b73a;
8'hfd : rvCrc[7] <= 32'hd0236bf0;
8'hfe : rvCrc[7] <= 32'h3cc10eae;
8'hff : rvCrc[7] <= 32'h6760d264;
endcase
case(iv_Input[071:064])
8'h00 : rvCrc[8] <= 32'h00000000;
8'h01 : rvCrc[8] <= 32'hf200aa66;
8'h02 : rvCrc[8] <= 32'he0c0497b;
8'h03 : rvCrc[8] <= 32'h12c0e31d;
8'h04 : rvCrc[8] <= 32'hc5418f41;
8'h05 : rvCrc[8] <= 32'h37412527;
8'h06 : rvCrc[8] <= 32'h2581c63a;
8'h07 : rvCrc[8] <= 32'hd7816c5c;
8'h08 : rvCrc[8] <= 32'h8e420335;
8'h09 : rvCrc[8] <= 32'h7c42a953;
8'h0a : rvCrc[8] <= 32'h6e824a4e;
8'h0b : rvCrc[8] <= 32'h9c82e028;
8'h0c : rvCrc[8] <= 32'h4b038c74;
8'h0d : rvCrc[8] <= 32'hb9032612;
8'h0e : rvCrc[8] <= 32'habc3c50f;
8'h0f : rvCrc[8] <= 32'h59c36f69;
8'h10 : rvCrc[8] <= 32'h18451bdd;
8'h11 : rvCrc[8] <= 32'hea45b1bb;
8'h12 : rvCrc[8] <= 32'hf88552a6;
8'h13 : rvCrc[8] <= 32'h0a85f8c0;
8'h14 : rvCrc[8] <= 32'hdd04949c;
8'h15 : rvCrc[8] <= 32'h2f043efa;
8'h16 : rvCrc[8] <= 32'h3dc4dde7;
8'h17 : rvCrc[8] <= 32'hcfc47781;
8'h18 : rvCrc[8] <= 32'h960718e8;
8'h19 : rvCrc[8] <= 32'h6407b28e;
8'h1a : rvCrc[8] <= 32'h76c75193;
8'h1b : rvCrc[8] <= 32'h84c7fbf5;
8'h1c : rvCrc[8] <= 32'h534697a9;
8'h1d : rvCrc[8] <= 32'ha1463dcf;
8'h1e : rvCrc[8] <= 32'hb386ded2;
8'h1f : rvCrc[8] <= 32'h418674b4;
8'h20 : rvCrc[8] <= 32'h308a37ba;
8'h21 : rvCrc[8] <= 32'hc28a9ddc;
8'h22 : rvCrc[8] <= 32'hd04a7ec1;
8'h23 : rvCrc[8] <= 32'h224ad4a7;
8'h24 : rvCrc[8] <= 32'hf5cbb8fb;
8'h25 : rvCrc[8] <= 32'h07cb129d;
8'h26 : rvCrc[8] <= 32'h150bf180;
8'h27 : rvCrc[8] <= 32'he70b5be6;
8'h28 : rvCrc[8] <= 32'hbec8348f;
8'h29 : rvCrc[8] <= 32'h4cc89ee9;
8'h2a : rvCrc[8] <= 32'h5e087df4;
8'h2b : rvCrc[8] <= 32'hac08d792;
8'h2c : rvCrc[8] <= 32'h7b89bbce;
8'h2d : rvCrc[8] <= 32'h898911a8;
8'h2e : rvCrc[8] <= 32'h9b49f2b5;
8'h2f : rvCrc[8] <= 32'h694958d3;
8'h30 : rvCrc[8] <= 32'h28cf2c67;
8'h31 : rvCrc[8] <= 32'hdacf8601;
8'h32 : rvCrc[8] <= 32'hc80f651c;
8'h33 : rvCrc[8] <= 32'h3a0fcf7a;
8'h34 : rvCrc[8] <= 32'hed8ea326;
8'h35 : rvCrc[8] <= 32'h1f8e0940;
8'h36 : rvCrc[8] <= 32'h0d4eea5d;
8'h37 : rvCrc[8] <= 32'hff4e403b;
8'h38 : rvCrc[8] <= 32'ha68d2f52;
8'h39 : rvCrc[8] <= 32'h548d8534;
8'h3a : rvCrc[8] <= 32'h464d6629;
8'h3b : rvCrc[8] <= 32'hb44dcc4f;
8'h3c : rvCrc[8] <= 32'h63cca013;
8'h3d : rvCrc[8] <= 32'h91cc0a75;
8'h3e : rvCrc[8] <= 32'h830ce968;
8'h3f : rvCrc[8] <= 32'h710c430e;
8'h40 : rvCrc[8] <= 32'h61146f74;
8'h41 : rvCrc[8] <= 32'h9314c512;
8'h42 : rvCrc[8] <= 32'h81d4260f;
8'h43 : rvCrc[8] <= 32'h73d48c69;
8'h44 : rvCrc[8] <= 32'ha455e035;
8'h45 : rvCrc[8] <= 32'h56554a53;
8'h46 : rvCrc[8] <= 32'h4495a94e;
8'h47 : rvCrc[8] <= 32'hb6950328;
8'h48 : rvCrc[8] <= 32'hef566c41;
8'h49 : rvCrc[8] <= 32'h1d56c627;
8'h4a : rvCrc[8] <= 32'h0f96253a;
8'h4b : rvCrc[8] <= 32'hfd968f5c;
8'h4c : rvCrc[8] <= 32'h2a17e300;
8'h4d : rvCrc[8] <= 32'hd8174966;
8'h4e : rvCrc[8] <= 32'hcad7aa7b;
8'h4f : rvCrc[8] <= 32'h38d7001d;
8'h50 : rvCrc[8] <= 32'h795174a9;
8'h51 : rvCrc[8] <= 32'h8b51decf;
8'h52 : rvCrc[8] <= 32'h99913dd2;
8'h53 : rvCrc[8] <= 32'h6b9197b4;
8'h54 : rvCrc[8] <= 32'hbc10fbe8;
8'h55 : rvCrc[8] <= 32'h4e10518e;
8'h56 : rvCrc[8] <= 32'h5cd0b293;
8'h57 : rvCrc[8] <= 32'haed018f5;
8'h58 : rvCrc[8] <= 32'hf713779c;
8'h59 : rvCrc[8] <= 32'h0513ddfa;
8'h5a : rvCrc[8] <= 32'h17d33ee7;
8'h5b : rvCrc[8] <= 32'he5d39481;
8'h5c : rvCrc[8] <= 32'h3252f8dd;
8'h5d : rvCrc[8] <= 32'hc05252bb;
8'h5e : rvCrc[8] <= 32'hd292b1a6;
8'h5f : rvCrc[8] <= 32'h20921bc0;
8'h60 : rvCrc[8] <= 32'h519e58ce;
8'h61 : rvCrc[8] <= 32'ha39ef2a8;
8'h62 : rvCrc[8] <= 32'hb15e11b5;
8'h63 : rvCrc[8] <= 32'h435ebbd3;
8'h64 : rvCrc[8] <= 32'h94dfd78f;
8'h65 : rvCrc[8] <= 32'h66df7de9;
8'h66 : rvCrc[8] <= 32'h741f9ef4;
8'h67 : rvCrc[8] <= 32'h861f3492;
8'h68 : rvCrc[8] <= 32'hdfdc5bfb;
8'h69 : rvCrc[8] <= 32'h2ddcf19d;
8'h6a : rvCrc[8] <= 32'h3f1c1280;
8'h6b : rvCrc[8] <= 32'hcd1cb8e6;
8'h6c : rvCrc[8] <= 32'h1a9dd4ba;
8'h6d : rvCrc[8] <= 32'he89d7edc;
8'h6e : rvCrc[8] <= 32'hfa5d9dc1;
8'h6f : rvCrc[8] <= 32'h085d37a7;
8'h70 : rvCrc[8] <= 32'h49db4313;
8'h71 : rvCrc[8] <= 32'hbbdbe975;
8'h72 : rvCrc[8] <= 32'ha91b0a68;
8'h73 : rvCrc[8] <= 32'h5b1ba00e;
8'h74 : rvCrc[8] <= 32'h8c9acc52;
8'h75 : rvCrc[8] <= 32'h7e9a6634;
8'h76 : rvCrc[8] <= 32'h6c5a8529;
8'h77 : rvCrc[8] <= 32'h9e5a2f4f;
8'h78 : rvCrc[8] <= 32'hc7994026;
8'h79 : rvCrc[8] <= 32'h3599ea40;
8'h7a : rvCrc[8] <= 32'h2759095d;
8'h7b : rvCrc[8] <= 32'hd559a33b;
8'h7c : rvCrc[8] <= 32'h02d8cf67;
8'h7d : rvCrc[8] <= 32'hf0d86501;
8'h7e : rvCrc[8] <= 32'he218861c;
8'h7f : rvCrc[8] <= 32'h10182c7a;
8'h80 : rvCrc[8] <= 32'hc228dee8;
8'h81 : rvCrc[8] <= 32'h3028748e;
8'h82 : rvCrc[8] <= 32'h22e89793;
8'h83 : rvCrc[8] <= 32'hd0e83df5;
8'h84 : rvCrc[8] <= 32'h076951a9;
8'h85 : rvCrc[8] <= 32'hf569fbcf;
8'h86 : rvCrc[8] <= 32'he7a918d2;
8'h87 : rvCrc[8] <= 32'h15a9b2b4;
8'h88 : rvCrc[8] <= 32'h4c6adddd;
8'h89 : rvCrc[8] <= 32'hbe6a77bb;
8'h8a : rvCrc[8] <= 32'hacaa94a6;
8'h8b : rvCrc[8] <= 32'h5eaa3ec0;
8'h8c : rvCrc[8] <= 32'h892b529c;
8'h8d : rvCrc[8] <= 32'h7b2bf8fa;
8'h8e : rvCrc[8] <= 32'h69eb1be7;
8'h8f : rvCrc[8] <= 32'h9bebb181;
8'h90 : rvCrc[8] <= 32'hda6dc535;
8'h91 : rvCrc[8] <= 32'h286d6f53;
8'h92 : rvCrc[8] <= 32'h3aad8c4e;
8'h93 : rvCrc[8] <= 32'hc8ad2628;
8'h94 : rvCrc[8] <= 32'h1f2c4a74;
8'h95 : rvCrc[8] <= 32'hed2ce012;
8'h96 : rvCrc[8] <= 32'hffec030f;
8'h97 : rvCrc[8] <= 32'h0deca969;
8'h98 : rvCrc[8] <= 32'h542fc600;
8'h99 : rvCrc[8] <= 32'ha62f6c66;
8'h9a : rvCrc[8] <= 32'hb4ef8f7b;
8'h9b : rvCrc[8] <= 32'h46ef251d;
8'h9c : rvCrc[8] <= 32'h916e4941;
8'h9d : rvCrc[8] <= 32'h636ee327;
8'h9e : rvCrc[8] <= 32'h71ae003a;
8'h9f : rvCrc[8] <= 32'h83aeaa5c;
8'ha0 : rvCrc[8] <= 32'hf2a2e952;
8'ha1 : rvCrc[8] <= 32'h00a24334;
8'ha2 : rvCrc[8] <= 32'h1262a029;
8'ha3 : rvCrc[8] <= 32'he0620a4f;
8'ha4 : rvCrc[8] <= 32'h37e36613;
8'ha5 : rvCrc[8] <= 32'hc5e3cc75;
8'ha6 : rvCrc[8] <= 32'hd7232f68;
8'ha7 : rvCrc[8] <= 32'h2523850e;
8'ha8 : rvCrc[8] <= 32'h7ce0ea67;
8'ha9 : rvCrc[8] <= 32'h8ee04001;
8'haa : rvCrc[8] <= 32'h9c20a31c;
8'hab : rvCrc[8] <= 32'h6e20097a;
8'hac : rvCrc[8] <= 32'hb9a16526;
8'had : rvCrc[8] <= 32'h4ba1cf40;
8'hae : rvCrc[8] <= 32'h59612c5d;
8'haf : rvCrc[8] <= 32'hab61863b;
8'hb0 : rvCrc[8] <= 32'heae7f28f;
8'hb1 : rvCrc[8] <= 32'h18e758e9;
8'hb2 : rvCrc[8] <= 32'h0a27bbf4;
8'hb3 : rvCrc[8] <= 32'hf8271192;
8'hb4 : rvCrc[8] <= 32'h2fa67dce;
8'hb5 : rvCrc[8] <= 32'hdda6d7a8;
8'hb6 : rvCrc[8] <= 32'hcf6634b5;
8'hb7 : rvCrc[8] <= 32'h3d669ed3;
8'hb8 : rvCrc[8] <= 32'h64a5f1ba;
8'hb9 : rvCrc[8] <= 32'h96a55bdc;
8'hba : rvCrc[8] <= 32'h8465b8c1;
8'hbb : rvCrc[8] <= 32'h766512a7;
8'hbc : rvCrc[8] <= 32'ha1e47efb;
8'hbd : rvCrc[8] <= 32'h53e4d49d;
8'hbe : rvCrc[8] <= 32'h41243780;
8'hbf : rvCrc[8] <= 32'hb3249de6;
8'hc0 : rvCrc[8] <= 32'ha33cb19c;
8'hc1 : rvCrc[8] <= 32'h513c1bfa;
8'hc2 : rvCrc[8] <= 32'h43fcf8e7;
8'hc3 : rvCrc[8] <= 32'hb1fc5281;
8'hc4 : rvCrc[8] <= 32'h667d3edd;
8'hc5 : rvCrc[8] <= 32'h947d94bb;
8'hc6 : rvCrc[8] <= 32'h86bd77a6;
8'hc7 : rvCrc[8] <= 32'h74bdddc0;
8'hc8 : rvCrc[8] <= 32'h2d7eb2a9;
8'hc9 : rvCrc[8] <= 32'hdf7e18cf;
8'hca : rvCrc[8] <= 32'hcdbefbd2;
8'hcb : rvCrc[8] <= 32'h3fbe51b4;
8'hcc : rvCrc[8] <= 32'he83f3de8;
8'hcd : rvCrc[8] <= 32'h1a3f978e;
8'hce : rvCrc[8] <= 32'h08ff7493;
8'hcf : rvCrc[8] <= 32'hfaffdef5;
8'hd0 : rvCrc[8] <= 32'hbb79aa41;
8'hd1 : rvCrc[8] <= 32'h49790027;
8'hd2 : rvCrc[8] <= 32'h5bb9e33a;
8'hd3 : rvCrc[8] <= 32'ha9b9495c;
8'hd4 : rvCrc[8] <= 32'h7e382500;
8'hd5 : rvCrc[8] <= 32'h8c388f66;
8'hd6 : rvCrc[8] <= 32'h9ef86c7b;
8'hd7 : rvCrc[8] <= 32'h6cf8c61d;
8'hd8 : rvCrc[8] <= 32'h353ba974;
8'hd9 : rvCrc[8] <= 32'hc73b0312;
8'hda : rvCrc[8] <= 32'hd5fbe00f;
8'hdb : rvCrc[8] <= 32'h27fb4a69;
8'hdc : rvCrc[8] <= 32'hf07a2635;
8'hdd : rvCrc[8] <= 32'h027a8c53;
8'hde : rvCrc[8] <= 32'h10ba6f4e;
8'hdf : rvCrc[8] <= 32'he2bac528;
8'he0 : rvCrc[8] <= 32'h93b68626;
8'he1 : rvCrc[8] <= 32'h61b62c40;
8'he2 : rvCrc[8] <= 32'h7376cf5d;
8'he3 : rvCrc[8] <= 32'h8176653b;
8'he4 : rvCrc[8] <= 32'h56f70967;
8'he5 : rvCrc[8] <= 32'ha4f7a301;
8'he6 : rvCrc[8] <= 32'hb637401c;
8'he7 : rvCrc[8] <= 32'h4437ea7a;
8'he8 : rvCrc[8] <= 32'h1df48513;
8'he9 : rvCrc[8] <= 32'heff42f75;
8'hea : rvCrc[8] <= 32'hfd34cc68;
8'heb : rvCrc[8] <= 32'h0f34660e;
8'hec : rvCrc[8] <= 32'hd8b50a52;
8'hed : rvCrc[8] <= 32'h2ab5a034;
8'hee : rvCrc[8] <= 32'h38754329;
8'hef : rvCrc[8] <= 32'hca75e94f;
8'hf0 : rvCrc[8] <= 32'h8bf39dfb;
8'hf1 : rvCrc[8] <= 32'h79f3379d;
8'hf2 : rvCrc[8] <= 32'h6b33d480;
8'hf3 : rvCrc[8] <= 32'h99337ee6;
8'hf4 : rvCrc[8] <= 32'h4eb212ba;
8'hf5 : rvCrc[8] <= 32'hbcb2b8dc;
8'hf6 : rvCrc[8] <= 32'hae725bc1;
8'hf7 : rvCrc[8] <= 32'h5c72f1a7;
8'hf8 : rvCrc[8] <= 32'h05b19ece;
8'hf9 : rvCrc[8] <= 32'hf7b134a8;
8'hfa : rvCrc[8] <= 32'he571d7b5;
8'hfb : rvCrc[8] <= 32'h17717dd3;
8'hfc : rvCrc[8] <= 32'hc0f0118f;
8'hfd : rvCrc[8] <= 32'h32f0bbe9;
8'hfe : rvCrc[8] <= 32'h203058f4;
8'hff : rvCrc[8] <= 32'hd230f292;
endcase
case(iv_Input[079:072])
8'h00 : rvCrc[9] <= 32'h00000000;
8'h01 : rvCrc[9] <= 32'h8090a067;
8'h02 : rvCrc[9] <= 32'h05e05d79;
8'h03 : rvCrc[9] <= 32'h8570fd1e;
8'h04 : rvCrc[9] <= 32'h0bc0baf2;
8'h05 : rvCrc[9] <= 32'h8b501a95;
8'h06 : rvCrc[9] <= 32'h0e20e78b;
8'h07 : rvCrc[9] <= 32'h8eb047ec;
8'h08 : rvCrc[9] <= 32'h178175e4;
8'h09 : rvCrc[9] <= 32'h9711d583;
8'h0a : rvCrc[9] <= 32'h1261289d;
8'h0b : rvCrc[9] <= 32'h92f188fa;
8'h0c : rvCrc[9] <= 32'h1c41cf16;
8'h0d : rvCrc[9] <= 32'h9cd16f71;
8'h0e : rvCrc[9] <= 32'h19a1926f;
8'h0f : rvCrc[9] <= 32'h99313208;
8'h10 : rvCrc[9] <= 32'h2f02ebc8;
8'h11 : rvCrc[9] <= 32'haf924baf;
8'h12 : rvCrc[9] <= 32'h2ae2b6b1;
8'h13 : rvCrc[9] <= 32'haa7216d6;
8'h14 : rvCrc[9] <= 32'h24c2513a;
8'h15 : rvCrc[9] <= 32'ha452f15d;
8'h16 : rvCrc[9] <= 32'h21220c43;
8'h17 : rvCrc[9] <= 32'ha1b2ac24;
8'h18 : rvCrc[9] <= 32'h38839e2c;
8'h19 : rvCrc[9] <= 32'hb8133e4b;
8'h1a : rvCrc[9] <= 32'h3d63c355;
8'h1b : rvCrc[9] <= 32'hbdf36332;
8'h1c : rvCrc[9] <= 32'h334324de;
8'h1d : rvCrc[9] <= 32'hb3d384b9;
8'h1e : rvCrc[9] <= 32'h36a379a7;
8'h1f : rvCrc[9] <= 32'hb633d9c0;
8'h20 : rvCrc[9] <= 32'h5e05d790;
8'h21 : rvCrc[9] <= 32'hde9577f7;
8'h22 : rvCrc[9] <= 32'h5be58ae9;
8'h23 : rvCrc[9] <= 32'hdb752a8e;
8'h24 : rvCrc[9] <= 32'h55c56d62;
8'h25 : rvCrc[9] <= 32'hd555cd05;
8'h26 : rvCrc[9] <= 32'h5025301b;
8'h27 : rvCrc[9] <= 32'hd0b5907c;
8'h28 : rvCrc[9] <= 32'h4984a274;
8'h29 : rvCrc[9] <= 32'hc9140213;
8'h2a : rvCrc[9] <= 32'h4c64ff0d;
8'h2b : rvCrc[9] <= 32'hccf45f6a;
8'h2c : rvCrc[9] <= 32'h42441886;
8'h2d : rvCrc[9] <= 32'hc2d4b8e1;
8'h2e : rvCrc[9] <= 32'h47a445ff;
8'h2f : rvCrc[9] <= 32'hc734e598;
8'h30 : rvCrc[9] <= 32'h71073c58;
8'h31 : rvCrc[9] <= 32'hf1979c3f;
8'h32 : rvCrc[9] <= 32'h74e76121;
8'h33 : rvCrc[9] <= 32'hf477c146;
8'h34 : rvCrc[9] <= 32'h7ac786aa;
8'h35 : rvCrc[9] <= 32'hfa5726cd;
8'h36 : rvCrc[9] <= 32'h7f27dbd3;
8'h37 : rvCrc[9] <= 32'hffb77bb4;
8'h38 : rvCrc[9] <= 32'h668649bc;
8'h39 : rvCrc[9] <= 32'he616e9db;
8'h3a : rvCrc[9] <= 32'h636614c5;
8'h3b : rvCrc[9] <= 32'he3f6b4a2;
8'h3c : rvCrc[9] <= 32'h6d46f34e;
8'h3d : rvCrc[9] <= 32'hedd65329;
8'h3e : rvCrc[9] <= 32'h68a6ae37;
8'h3f : rvCrc[9] <= 32'he8360e50;
8'h40 : rvCrc[9] <= 32'hbc0baf20;
8'h41 : rvCrc[9] <= 32'h3c9b0f47;
8'h42 : rvCrc[9] <= 32'hb9ebf259;
8'h43 : rvCrc[9] <= 32'h397b523e;
8'h44 : rvCrc[9] <= 32'hb7cb15d2;
8'h45 : rvCrc[9] <= 32'h375bb5b5;
8'h46 : rvCrc[9] <= 32'hb22b48ab;
8'h47 : rvCrc[9] <= 32'h32bbe8cc;
8'h48 : rvCrc[9] <= 32'hab8adac4;
8'h49 : rvCrc[9] <= 32'h2b1a7aa3;
8'h4a : rvCrc[9] <= 32'hae6a87bd;
8'h4b : rvCrc[9] <= 32'h2efa27da;
8'h4c : rvCrc[9] <= 32'ha04a6036;
8'h4d : rvCrc[9] <= 32'h20dac051;
8'h4e : rvCrc[9] <= 32'ha5aa3d4f;
8'h4f : rvCrc[9] <= 32'h253a9d28;
8'h50 : rvCrc[9] <= 32'h930944e8;
8'h51 : rvCrc[9] <= 32'h1399e48f;
8'h52 : rvCrc[9] <= 32'h96e91991;
8'h53 : rvCrc[9] <= 32'h1679b9f6;
8'h54 : rvCrc[9] <= 32'h98c9fe1a;
8'h55 : rvCrc[9] <= 32'h18595e7d;
8'h56 : rvCrc[9] <= 32'h9d29a363;
8'h57 : rvCrc[9] <= 32'h1db90304;
8'h58 : rvCrc[9] <= 32'h8488310c;
8'h59 : rvCrc[9] <= 32'h0418916b;
8'h5a : rvCrc[9] <= 32'h81686c75;
8'h5b : rvCrc[9] <= 32'h01f8cc12;
8'h5c : rvCrc[9] <= 32'h8f488bfe;
8'h5d : rvCrc[9] <= 32'h0fd82b99;
8'h5e : rvCrc[9] <= 32'h8aa8d687;
8'h5f : rvCrc[9] <= 32'h0a3876e0;
8'h60 : rvCrc[9] <= 32'he20e78b0;
8'h61 : rvCrc[9] <= 32'h629ed8d7;
8'h62 : rvCrc[9] <= 32'he7ee25c9;
8'h63 : rvCrc[9] <= 32'h677e85ae;
8'h64 : rvCrc[9] <= 32'he9cec242;
8'h65 : rvCrc[9] <= 32'h695e6225;
8'h66 : rvCrc[9] <= 32'hec2e9f3b;
8'h67 : rvCrc[9] <= 32'h6cbe3f5c;
8'h68 : rvCrc[9] <= 32'hf58f0d54;
8'h69 : rvCrc[9] <= 32'h751fad33;
8'h6a : rvCrc[9] <= 32'hf06f502d;
8'h6b : rvCrc[9] <= 32'h70fff04a;
8'h6c : rvCrc[9] <= 32'hfe4fb7a6;
8'h6d : rvCrc[9] <= 32'h7edf17c1;
8'h6e : rvCrc[9] <= 32'hfbafeadf;
8'h6f : rvCrc[9] <= 32'h7b3f4ab8;
8'h70 : rvCrc[9] <= 32'hcd0c9378;
8'h71 : rvCrc[9] <= 32'h4d9c331f;
8'h72 : rvCrc[9] <= 32'hc8ecce01;
8'h73 : rvCrc[9] <= 32'h487c6e66;
8'h74 : rvCrc[9] <= 32'hc6cc298a;
8'h75 : rvCrc[9] <= 32'h465c89ed;
8'h76 : rvCrc[9] <= 32'hc32c74f3;
8'h77 : rvCrc[9] <= 32'h43bcd494;
8'h78 : rvCrc[9] <= 32'hda8de69c;
8'h79 : rvCrc[9] <= 32'h5a1d46fb;
8'h7a : rvCrc[9] <= 32'hdf6dbbe5;
8'h7b : rvCrc[9] <= 32'h5ffd1b82;
8'h7c : rvCrc[9] <= 32'hd14d5c6e;
8'h7d : rvCrc[9] <= 32'h51ddfc09;
8'h7e : rvCrc[9] <= 32'hd4ad0117;
8'h7f : rvCrc[9] <= 32'h543da170;
8'h80 : rvCrc[9] <= 32'h7cd643f7;
8'h81 : rvCrc[9] <= 32'hfc46e390;
8'h82 : rvCrc[9] <= 32'h79361e8e;
8'h83 : rvCrc[9] <= 32'hf9a6bee9;
8'h84 : rvCrc[9] <= 32'h7716f905;
8'h85 : rvCrc[9] <= 32'hf7865962;
8'h86 : rvCrc[9] <= 32'h72f6a47c;
8'h87 : rvCrc[9] <= 32'hf266041b;
8'h88 : rvCrc[9] <= 32'h6b573613;
8'h89 : rvCrc[9] <= 32'hebc79674;
8'h8a : rvCrc[9] <= 32'h6eb76b6a;
8'h8b : rvCrc[9] <= 32'hee27cb0d;
8'h8c : rvCrc[9] <= 32'h60978ce1;
8'h8d : rvCrc[9] <= 32'he0072c86;
8'h8e : rvCrc[9] <= 32'h6577d198;
8'h8f : rvCrc[9] <= 32'he5e771ff;
8'h90 : rvCrc[9] <= 32'h53d4a83f;
8'h91 : rvCrc[9] <= 32'hd3440858;
8'h92 : rvCrc[9] <= 32'h5634f546;
8'h93 : rvCrc[9] <= 32'hd6a45521;
8'h94 : rvCrc[9] <= 32'h581412cd;
8'h95 : rvCrc[9] <= 32'hd884b2aa;
8'h96 : rvCrc[9] <= 32'h5df44fb4;
8'h97 : rvCrc[9] <= 32'hdd64efd3;
8'h98 : rvCrc[9] <= 32'h4455dddb;
8'h99 : rvCrc[9] <= 32'hc4c57dbc;
8'h9a : rvCrc[9] <= 32'h41b580a2;
8'h9b : rvCrc[9] <= 32'hc12520c5;
8'h9c : rvCrc[9] <= 32'h4f956729;
8'h9d : rvCrc[9] <= 32'hcf05c74e;
8'h9e : rvCrc[9] <= 32'h4a753a50;
8'h9f : rvCrc[9] <= 32'hcae59a37;
8'ha0 : rvCrc[9] <= 32'h22d39467;
8'ha1 : rvCrc[9] <= 32'ha2433400;
8'ha2 : rvCrc[9] <= 32'h2733c91e;
8'ha3 : rvCrc[9] <= 32'ha7a36979;
8'ha4 : rvCrc[9] <= 32'h29132e95;
8'ha5 : rvCrc[9] <= 32'ha9838ef2;
8'ha6 : rvCrc[9] <= 32'h2cf373ec;
8'ha7 : rvCrc[9] <= 32'hac63d38b;
8'ha8 : rvCrc[9] <= 32'h3552e183;
8'ha9 : rvCrc[9] <= 32'hb5c241e4;
8'haa : rvCrc[9] <= 32'h30b2bcfa;
8'hab : rvCrc[9] <= 32'hb0221c9d;
8'hac : rvCrc[9] <= 32'h3e925b71;
8'had : rvCrc[9] <= 32'hbe02fb16;
8'hae : rvCrc[9] <= 32'h3b720608;
8'haf : rvCrc[9] <= 32'hbbe2a66f;
8'hb0 : rvCrc[9] <= 32'h0dd17faf;
8'hb1 : rvCrc[9] <= 32'h8d41dfc8;
8'hb2 : rvCrc[9] <= 32'h083122d6;
8'hb3 : rvCrc[9] <= 32'h88a182b1;
8'hb4 : rvCrc[9] <= 32'h0611c55d;
8'hb5 : rvCrc[9] <= 32'h8681653a;
8'hb6 : rvCrc[9] <= 32'h03f19824;
8'hb7 : rvCrc[9] <= 32'h83613843;
8'hb8 : rvCrc[9] <= 32'h1a500a4b;
8'hb9 : rvCrc[9] <= 32'h9ac0aa2c;
8'hba : rvCrc[9] <= 32'h1fb05732;
8'hbb : rvCrc[9] <= 32'h9f20f755;
8'hbc : rvCrc[9] <= 32'h1190b0b9;
8'hbd : rvCrc[9] <= 32'h910010de;
8'hbe : rvCrc[9] <= 32'h1470edc0;
8'hbf : rvCrc[9] <= 32'h94e04da7;
8'hc0 : rvCrc[9] <= 32'hc0ddecd7;
8'hc1 : rvCrc[9] <= 32'h404d4cb0;
8'hc2 : rvCrc[9] <= 32'hc53db1ae;
8'hc3 : rvCrc[9] <= 32'h45ad11c9;
8'hc4 : rvCrc[9] <= 32'hcb1d5625;
8'hc5 : rvCrc[9] <= 32'h4b8df642;
8'hc6 : rvCrc[9] <= 32'hcefd0b5c;
8'hc7 : rvCrc[9] <= 32'h4e6dab3b;
8'hc8 : rvCrc[9] <= 32'hd75c9933;
8'hc9 : rvCrc[9] <= 32'h57cc3954;
8'hca : rvCrc[9] <= 32'hd2bcc44a;
8'hcb : rvCrc[9] <= 32'h522c642d;
8'hcc : rvCrc[9] <= 32'hdc9c23c1;
8'hcd : rvCrc[9] <= 32'h5c0c83a6;
8'hce : rvCrc[9] <= 32'hd97c7eb8;
8'hcf : rvCrc[9] <= 32'h59ecdedf;
8'hd0 : rvCrc[9] <= 32'hefdf071f;
8'hd1 : rvCrc[9] <= 32'h6f4fa778;
8'hd2 : rvCrc[9] <= 32'hea3f5a66;
8'hd3 : rvCrc[9] <= 32'h6aaffa01;
8'hd4 : rvCrc[9] <= 32'he41fbded;
8'hd5 : rvCrc[9] <= 32'h648f1d8a;
8'hd6 : rvCrc[9] <= 32'he1ffe094;
8'hd7 : rvCrc[9] <= 32'h616f40f3;
8'hd8 : rvCrc[9] <= 32'hf85e72fb;
8'hd9 : rvCrc[9] <= 32'h78ced29c;
8'hda : rvCrc[9] <= 32'hfdbe2f82;
8'hdb : rvCrc[9] <= 32'h7d2e8fe5;
8'hdc : rvCrc[9] <= 32'hf39ec809;
8'hdd : rvCrc[9] <= 32'h730e686e;
8'hde : rvCrc[9] <= 32'hf67e9570;
8'hdf : rvCrc[9] <= 32'h76ee3517;
8'he0 : rvCrc[9] <= 32'h9ed83b47;
8'he1 : rvCrc[9] <= 32'h1e489b20;
8'he2 : rvCrc[9] <= 32'h9b38663e;
8'he3 : rvCrc[9] <= 32'h1ba8c659;
8'he4 : rvCrc[9] <= 32'h951881b5;
8'he5 : rvCrc[9] <= 32'h158821d2;
8'he6 : rvCrc[9] <= 32'h90f8dccc;
8'he7 : rvCrc[9] <= 32'h10687cab;
8'he8 : rvCrc[9] <= 32'h89594ea3;
8'he9 : rvCrc[9] <= 32'h09c9eec4;
8'hea : rvCrc[9] <= 32'h8cb913da;
8'heb : rvCrc[9] <= 32'h0c29b3bd;
8'hec : rvCrc[9] <= 32'h8299f451;
8'hed : rvCrc[9] <= 32'h02095436;
8'hee : rvCrc[9] <= 32'h8779a928;
8'hef : rvCrc[9] <= 32'h07e9094f;
8'hf0 : rvCrc[9] <= 32'hb1dad08f;
8'hf1 : rvCrc[9] <= 32'h314a70e8;
8'hf2 : rvCrc[9] <= 32'hb43a8df6;
8'hf3 : rvCrc[9] <= 32'h34aa2d91;
8'hf4 : rvCrc[9] <= 32'hba1a6a7d;
8'hf5 : rvCrc[9] <= 32'h3a8aca1a;
8'hf6 : rvCrc[9] <= 32'hbffa3704;
8'hf7 : rvCrc[9] <= 32'h3f6a9763;
8'hf8 : rvCrc[9] <= 32'ha65ba56b;
8'hf9 : rvCrc[9] <= 32'h26cb050c;
8'hfa : rvCrc[9] <= 32'ha3bbf812;
8'hfb : rvCrc[9] <= 32'h232b5875;
8'hfc : rvCrc[9] <= 32'had9b1f99;
8'hfd : rvCrc[9] <= 32'h2d0bbffe;
8'hfe : rvCrc[9] <= 32'ha87b42e0;
8'hff : rvCrc[9] <= 32'h28ebe287;
endcase
case(iv_Input[087:080])
8'h00 : rvCrc[10] <= 32'h00000000;
8'h01 : rvCrc[10] <= 32'hf9ac87ee;
8'h02 : rvCrc[10] <= 32'hf798126b;
8'h03 : rvCrc[10] <= 32'h0e349585;
8'h04 : rvCrc[10] <= 32'hebf13961;
8'h05 : rvCrc[10] <= 32'h125dbe8f;
8'h06 : rvCrc[10] <= 32'h1c692b0a;
8'h07 : rvCrc[10] <= 32'he5c5ace4;
8'h08 : rvCrc[10] <= 32'hd3236f75;
8'h09 : rvCrc[10] <= 32'h2a8fe89b;
8'h0a : rvCrc[10] <= 32'h24bb7d1e;
8'h0b : rvCrc[10] <= 32'hdd17faf0;
8'h0c : rvCrc[10] <= 32'h38d25614;
8'h0d : rvCrc[10] <= 32'hc17ed1fa;
8'h0e : rvCrc[10] <= 32'hcf4a447f;
8'h0f : rvCrc[10] <= 32'h36e6c391;
8'h10 : rvCrc[10] <= 32'ha287c35d;
8'h11 : rvCrc[10] <= 32'h5b2b44b3;
8'h12 : rvCrc[10] <= 32'h551fd136;
8'h13 : rvCrc[10] <= 32'hacb356d8;
8'h14 : rvCrc[10] <= 32'h4976fa3c;
8'h15 : rvCrc[10] <= 32'hb0da7dd2;
8'h16 : rvCrc[10] <= 32'hbeeee857;
8'h17 : rvCrc[10] <= 32'h47426fb9;
8'h18 : rvCrc[10] <= 32'h71a4ac28;
8'h19 : rvCrc[10] <= 32'h88082bc6;
8'h1a : rvCrc[10] <= 32'h863cbe43;
8'h1b : rvCrc[10] <= 32'h7f9039ad;
8'h1c : rvCrc[10] <= 32'h9a559549;
8'h1d : rvCrc[10] <= 32'h63f912a7;
8'h1e : rvCrc[10] <= 32'h6dcd8722;
8'h1f : rvCrc[10] <= 32'h946100cc;
8'h20 : rvCrc[10] <= 32'h41ce9b0d;
8'h21 : rvCrc[10] <= 32'hb8621ce3;
8'h22 : rvCrc[10] <= 32'hb6568966;
8'h23 : rvCrc[10] <= 32'h4ffa0e88;
8'h24 : rvCrc[10] <= 32'haa3fa26c;
8'h25 : rvCrc[10] <= 32'h53932582;
8'h26 : rvCrc[10] <= 32'h5da7b007;
8'h27 : rvCrc[10] <= 32'ha40b37e9;
8'h28 : rvCrc[10] <= 32'h92edf478;
8'h29 : rvCrc[10] <= 32'h6b417396;
8'h2a : rvCrc[10] <= 32'h6575e613;
8'h2b : rvCrc[10] <= 32'h9cd961fd;
8'h2c : rvCrc[10] <= 32'h791ccd19;
8'h2d : rvCrc[10] <= 32'h80b04af7;
8'h2e : rvCrc[10] <= 32'h8e84df72;
8'h2f : rvCrc[10] <= 32'h7728589c;
8'h30 : rvCrc[10] <= 32'he3495850;
8'h31 : rvCrc[10] <= 32'h1ae5dfbe;
8'h32 : rvCrc[10] <= 32'h14d14a3b;
8'h33 : rvCrc[10] <= 32'hed7dcdd5;
8'h34 : rvCrc[10] <= 32'h08b86131;
8'h35 : rvCrc[10] <= 32'hf114e6df;
8'h36 : rvCrc[10] <= 32'hff20735a;
8'h37 : rvCrc[10] <= 32'h068cf4b4;
8'h38 : rvCrc[10] <= 32'h306a3725;
8'h39 : rvCrc[10] <= 32'hc9c6b0cb;
8'h3a : rvCrc[10] <= 32'hc7f2254e;
8'h3b : rvCrc[10] <= 32'h3e5ea2a0;
8'h3c : rvCrc[10] <= 32'hdb9b0e44;
8'h3d : rvCrc[10] <= 32'h223789aa;
8'h3e : rvCrc[10] <= 32'h2c031c2f;
8'h3f : rvCrc[10] <= 32'hd5af9bc1;
8'h40 : rvCrc[10] <= 32'h839d361a;
8'h41 : rvCrc[10] <= 32'h7a31b1f4;
8'h42 : rvCrc[10] <= 32'h74052471;
8'h43 : rvCrc[10] <= 32'h8da9a39f;
8'h44 : rvCrc[10] <= 32'h686c0f7b;
8'h45 : rvCrc[10] <= 32'h91c08895;
8'h46 : rvCrc[10] <= 32'h9ff41d10;
8'h47 : rvCrc[10] <= 32'h66589afe;
8'h48 : rvCrc[10] <= 32'h50be596f;
8'h49 : rvCrc[10] <= 32'ha912de81;
8'h4a : rvCrc[10] <= 32'ha7264b04;
8'h4b : rvCrc[10] <= 32'h5e8accea;
8'h4c : rvCrc[10] <= 32'hbb4f600e;
8'h4d : rvCrc[10] <= 32'h42e3e7e0;
8'h4e : rvCrc[10] <= 32'h4cd77265;
8'h4f : rvCrc[10] <= 32'hb57bf58b;
8'h50 : rvCrc[10] <= 32'h211af547;
8'h51 : rvCrc[10] <= 32'hd8b672a9;
8'h52 : rvCrc[10] <= 32'hd682e72c;
8'h53 : rvCrc[10] <= 32'h2f2e60c2;
8'h54 : rvCrc[10] <= 32'hcaebcc26;
8'h55 : rvCrc[10] <= 32'h33474bc8;
8'h56 : rvCrc[10] <= 32'h3d73de4d;
8'h57 : rvCrc[10] <= 32'hc4df59a3;
8'h58 : rvCrc[10] <= 32'hf2399a32;
8'h59 : rvCrc[10] <= 32'h0b951ddc;
8'h5a : rvCrc[10] <= 32'h05a18859;
8'h5b : rvCrc[10] <= 32'hfc0d0fb7;
8'h5c : rvCrc[10] <= 32'h19c8a353;
8'h5d : rvCrc[10] <= 32'he06424bd;
8'h5e : rvCrc[10] <= 32'hee50b138;
8'h5f : rvCrc[10] <= 32'h17fc36d6;
8'h60 : rvCrc[10] <= 32'hc253ad17;
8'h61 : rvCrc[10] <= 32'h3bff2af9;
8'h62 : rvCrc[10] <= 32'h35cbbf7c;
8'h63 : rvCrc[10] <= 32'hcc673892;
8'h64 : rvCrc[10] <= 32'h29a29476;
8'h65 : rvCrc[10] <= 32'hd00e1398;
8'h66 : rvCrc[10] <= 32'hde3a861d;
8'h67 : rvCrc[10] <= 32'h279601f3;
8'h68 : rvCrc[10] <= 32'h1170c262;
8'h69 : rvCrc[10] <= 32'he8dc458c;
8'h6a : rvCrc[10] <= 32'he6e8d009;
8'h6b : rvCrc[10] <= 32'h1f4457e7;
8'h6c : rvCrc[10] <= 32'hfa81fb03;
8'h6d : rvCrc[10] <= 32'h032d7ced;
8'h6e : rvCrc[10] <= 32'h0d19e968;
8'h6f : rvCrc[10] <= 32'hf4b56e86;
8'h70 : rvCrc[10] <= 32'h60d46e4a;
8'h71 : rvCrc[10] <= 32'h9978e9a4;
8'h72 : rvCrc[10] <= 32'h974c7c21;
8'h73 : rvCrc[10] <= 32'h6ee0fbcf;
8'h74 : rvCrc[10] <= 32'h8b25572b;
8'h75 : rvCrc[10] <= 32'h7289d0c5;
8'h76 : rvCrc[10] <= 32'h7cbd4540;
8'h77 : rvCrc[10] <= 32'h8511c2ae;
8'h78 : rvCrc[10] <= 32'hb3f7013f;
8'h79 : rvCrc[10] <= 32'h4a5b86d1;
8'h7a : rvCrc[10] <= 32'h446f1354;
8'h7b : rvCrc[10] <= 32'hbdc394ba;
8'h7c : rvCrc[10] <= 32'h5806385e;
8'h7d : rvCrc[10] <= 32'ha1aabfb0;
8'h7e : rvCrc[10] <= 32'haf9e2a35;
8'h7f : rvCrc[10] <= 32'h5632addb;
8'h80 : rvCrc[10] <= 32'h03fb7183;
8'h81 : rvCrc[10] <= 32'hfa57f66d;
8'h82 : rvCrc[10] <= 32'hf46363e8;
8'h83 : rvCrc[10] <= 32'h0dcfe406;
8'h84 : rvCrc[10] <= 32'he80a48e2;
8'h85 : rvCrc[10] <= 32'h11a6cf0c;
8'h86 : rvCrc[10] <= 32'h1f925a89;
8'h87 : rvCrc[10] <= 32'he63edd67;
8'h88 : rvCrc[10] <= 32'hd0d81ef6;
8'h89 : rvCrc[10] <= 32'h29749918;
8'h8a : rvCrc[10] <= 32'h27400c9d;
8'h8b : rvCrc[10] <= 32'hdeec8b73;
8'h8c : rvCrc[10] <= 32'h3b292797;
8'h8d : rvCrc[10] <= 32'hc285a079;
8'h8e : rvCrc[10] <= 32'hccb135fc;
8'h8f : rvCrc[10] <= 32'h351db212;
8'h90 : rvCrc[10] <= 32'ha17cb2de;
8'h91 : rvCrc[10] <= 32'h58d03530;
8'h92 : rvCrc[10] <= 32'h56e4a0b5;
8'h93 : rvCrc[10] <= 32'haf48275b;
8'h94 : rvCrc[10] <= 32'h4a8d8bbf;
8'h95 : rvCrc[10] <= 32'hb3210c51;
8'h96 : rvCrc[10] <= 32'hbd1599d4;
8'h97 : rvCrc[10] <= 32'h44b91e3a;
8'h98 : rvCrc[10] <= 32'h725fddab;
8'h99 : rvCrc[10] <= 32'h8bf35a45;
8'h9a : rvCrc[10] <= 32'h85c7cfc0;
8'h9b : rvCrc[10] <= 32'h7c6b482e;
8'h9c : rvCrc[10] <= 32'h99aee4ca;
8'h9d : rvCrc[10] <= 32'h60026324;
8'h9e : rvCrc[10] <= 32'h6e36f6a1;
8'h9f : rvCrc[10] <= 32'h979a714f;
8'ha0 : rvCrc[10] <= 32'h4235ea8e;
8'ha1 : rvCrc[10] <= 32'hbb996d60;
8'ha2 : rvCrc[10] <= 32'hb5adf8e5;
8'ha3 : rvCrc[10] <= 32'h4c017f0b;
8'ha4 : rvCrc[10] <= 32'ha9c4d3ef;
8'ha5 : rvCrc[10] <= 32'h50685401;
8'ha6 : rvCrc[10] <= 32'h5e5cc184;
8'ha7 : rvCrc[10] <= 32'ha7f0466a;
8'ha8 : rvCrc[10] <= 32'h911685fb;
8'ha9 : rvCrc[10] <= 32'h68ba0215;
8'haa : rvCrc[10] <= 32'h668e9790;
8'hab : rvCrc[10] <= 32'h9f22107e;
8'hac : rvCrc[10] <= 32'h7ae7bc9a;
8'had : rvCrc[10] <= 32'h834b3b74;
8'hae : rvCrc[10] <= 32'h8d7faef1;
8'haf : rvCrc[10] <= 32'h74d3291f;
8'hb0 : rvCrc[10] <= 32'he0b229d3;
8'hb1 : rvCrc[10] <= 32'h191eae3d;
8'hb2 : rvCrc[10] <= 32'h172a3bb8;
8'hb3 : rvCrc[10] <= 32'hee86bc56;
8'hb4 : rvCrc[10] <= 32'h0b4310b2;
8'hb5 : rvCrc[10] <= 32'hf2ef975c;
8'hb6 : rvCrc[10] <= 32'hfcdb02d9;
8'hb7 : rvCrc[10] <= 32'h05778537;
8'hb8 : rvCrc[10] <= 32'h339146a6;
8'hb9 : rvCrc[10] <= 32'hca3dc148;
8'hba : rvCrc[10] <= 32'hc40954cd;
8'hbb : rvCrc[10] <= 32'h3da5d323;
8'hbc : rvCrc[10] <= 32'hd8607fc7;
8'hbd : rvCrc[10] <= 32'h21ccf829;
8'hbe : rvCrc[10] <= 32'h2ff86dac;
8'hbf : rvCrc[10] <= 32'hd654ea42;
8'hc0 : rvCrc[10] <= 32'h80664799;
8'hc1 : rvCrc[10] <= 32'h79cac077;
8'hc2 : rvCrc[10] <= 32'h77fe55f2;
8'hc3 : rvCrc[10] <= 32'h8e52d21c;
8'hc4 : rvCrc[10] <= 32'h6b977ef8;
8'hc5 : rvCrc[10] <= 32'h923bf916;
8'hc6 : rvCrc[10] <= 32'h9c0f6c93;
8'hc7 : rvCrc[10] <= 32'h65a3eb7d;
8'hc8 : rvCrc[10] <= 32'h534528ec;
8'hc9 : rvCrc[10] <= 32'haae9af02;
8'hca : rvCrc[10] <= 32'ha4dd3a87;
8'hcb : rvCrc[10] <= 32'h5d71bd69;
8'hcc : rvCrc[10] <= 32'hb8b4118d;
8'hcd : rvCrc[10] <= 32'h41189663;
8'hce : rvCrc[10] <= 32'h4f2c03e6;
8'hcf : rvCrc[10] <= 32'hb6808408;
8'hd0 : rvCrc[10] <= 32'h22e184c4;
8'hd1 : rvCrc[10] <= 32'hdb4d032a;
8'hd2 : rvCrc[10] <= 32'hd57996af;
8'hd3 : rvCrc[10] <= 32'h2cd51141;
8'hd4 : rvCrc[10] <= 32'hc910bda5;
8'hd5 : rvCrc[10] <= 32'h30bc3a4b;
8'hd6 : rvCrc[10] <= 32'h3e88afce;
8'hd7 : rvCrc[10] <= 32'hc7242820;
8'hd8 : rvCrc[10] <= 32'hf1c2ebb1;
8'hd9 : rvCrc[10] <= 32'h086e6c5f;
8'hda : rvCrc[10] <= 32'h065af9da;
8'hdb : rvCrc[10] <= 32'hfff67e34;
8'hdc : rvCrc[10] <= 32'h1a33d2d0;
8'hdd : rvCrc[10] <= 32'he39f553e;
8'hde : rvCrc[10] <= 32'hedabc0bb;
8'hdf : rvCrc[10] <= 32'h14074755;
8'he0 : rvCrc[10] <= 32'hc1a8dc94;
8'he1 : rvCrc[10] <= 32'h38045b7a;
8'he2 : rvCrc[10] <= 32'h3630ceff;
8'he3 : rvCrc[10] <= 32'hcf9c4911;
8'he4 : rvCrc[10] <= 32'h2a59e5f5;
8'he5 : rvCrc[10] <= 32'hd3f5621b;
8'he6 : rvCrc[10] <= 32'hddc1f79e;
8'he7 : rvCrc[10] <= 32'h246d7070;
8'he8 : rvCrc[10] <= 32'h128bb3e1;
8'he9 : rvCrc[10] <= 32'heb27340f;
8'hea : rvCrc[10] <= 32'he513a18a;
8'heb : rvCrc[10] <= 32'h1cbf2664;
8'hec : rvCrc[10] <= 32'hf97a8a80;
8'hed : rvCrc[10] <= 32'h00d60d6e;
8'hee : rvCrc[10] <= 32'h0ee298eb;
8'hef : rvCrc[10] <= 32'hf74e1f05;
8'hf0 : rvCrc[10] <= 32'h632f1fc9;
8'hf1 : rvCrc[10] <= 32'h9a839827;
8'hf2 : rvCrc[10] <= 32'h94b70da2;
8'hf3 : rvCrc[10] <= 32'h6d1b8a4c;
8'hf4 : rvCrc[10] <= 32'h88de26a8;
8'hf5 : rvCrc[10] <= 32'h7172a146;
8'hf6 : rvCrc[10] <= 32'h7f4634c3;
8'hf7 : rvCrc[10] <= 32'h86eab32d;
8'hf8 : rvCrc[10] <= 32'hb00c70bc;
8'hf9 : rvCrc[10] <= 32'h49a0f752;
8'hfa : rvCrc[10] <= 32'h479462d7;
8'hfb : rvCrc[10] <= 32'hbe38e539;
8'hfc : rvCrc[10] <= 32'h5bfd49dd;
8'hfd : rvCrc[10] <= 32'ha251ce33;
8'hfe : rvCrc[10] <= 32'hac655bb6;
8'hff : rvCrc[10] <= 32'h55c9dc58;
endcase
case(iv_Input[095:088])
8'h00 : rvCrc[11] <= 32'h00000000;
8'h01 : rvCrc[11] <= 32'h07f6e306;
8'h02 : rvCrc[11] <= 32'h0fedc60c;
8'h03 : rvCrc[11] <= 32'h081b250a;
8'h04 : rvCrc[11] <= 32'h1fdb8c18;
8'h05 : rvCrc[11] <= 32'h182d6f1e;
8'h06 : rvCrc[11] <= 32'h10364a14;
8'h07 : rvCrc[11] <= 32'h17c0a912;
8'h08 : rvCrc[11] <= 32'h3fb71830;
8'h09 : rvCrc[11] <= 32'h3841fb36;
8'h0a : rvCrc[11] <= 32'h305ade3c;
8'h0b : rvCrc[11] <= 32'h37ac3d3a;
8'h0c : rvCrc[11] <= 32'h206c9428;
8'h0d : rvCrc[11] <= 32'h279a772e;
8'h0e : rvCrc[11] <= 32'h2f815224;
8'h0f : rvCrc[11] <= 32'h2877b122;
8'h10 : rvCrc[11] <= 32'h7f6e3060;
8'h11 : rvCrc[11] <= 32'h7898d366;
8'h12 : rvCrc[11] <= 32'h7083f66c;
8'h13 : rvCrc[11] <= 32'h7775156a;
8'h14 : rvCrc[11] <= 32'h60b5bc78;
8'h15 : rvCrc[11] <= 32'h67435f7e;
8'h16 : rvCrc[11] <= 32'h6f587a74;
8'h17 : rvCrc[11] <= 32'h68ae9972;
8'h18 : rvCrc[11] <= 32'h40d92850;
8'h19 : rvCrc[11] <= 32'h472fcb56;
8'h1a : rvCrc[11] <= 32'h4f34ee5c;
8'h1b : rvCrc[11] <= 32'h48c20d5a;
8'h1c : rvCrc[11] <= 32'h5f02a448;
8'h1d : rvCrc[11] <= 32'h58f4474e;
8'h1e : rvCrc[11] <= 32'h50ef6244;
8'h1f : rvCrc[11] <= 32'h57198142;
8'h20 : rvCrc[11] <= 32'hfedc60c0;
8'h21 : rvCrc[11] <= 32'hf92a83c6;
8'h22 : rvCrc[11] <= 32'hf131a6cc;
8'h23 : rvCrc[11] <= 32'hf6c745ca;
8'h24 : rvCrc[11] <= 32'he107ecd8;
8'h25 : rvCrc[11] <= 32'he6f10fde;
8'h26 : rvCrc[11] <= 32'heeea2ad4;
8'h27 : rvCrc[11] <= 32'he91cc9d2;
8'h28 : rvCrc[11] <= 32'hc16b78f0;
8'h29 : rvCrc[11] <= 32'hc69d9bf6;
8'h2a : rvCrc[11] <= 32'hce86befc;
8'h2b : rvCrc[11] <= 32'hc9705dfa;
8'h2c : rvCrc[11] <= 32'hdeb0f4e8;
8'h2d : rvCrc[11] <= 32'hd94617ee;
8'h2e : rvCrc[11] <= 32'hd15d32e4;
8'h2f : rvCrc[11] <= 32'hd6abd1e2;
8'h30 : rvCrc[11] <= 32'h81b250a0;
8'h31 : rvCrc[11] <= 32'h8644b3a6;
8'h32 : rvCrc[11] <= 32'h8e5f96ac;
8'h33 : rvCrc[11] <= 32'h89a975aa;
8'h34 : rvCrc[11] <= 32'h9e69dcb8;
8'h35 : rvCrc[11] <= 32'h999f3fbe;
8'h36 : rvCrc[11] <= 32'h91841ab4;
8'h37 : rvCrc[11] <= 32'h9672f9b2;
8'h38 : rvCrc[11] <= 32'hbe054890;
8'h39 : rvCrc[11] <= 32'hb9f3ab96;
8'h3a : rvCrc[11] <= 32'hb1e88e9c;
8'h3b : rvCrc[11] <= 32'hb61e6d9a;
8'h3c : rvCrc[11] <= 32'ha1dec488;
8'h3d : rvCrc[11] <= 32'ha628278e;
8'h3e : rvCrc[11] <= 32'hae330284;
8'h3f : rvCrc[11] <= 32'ha9c5e182;
8'h40 : rvCrc[11] <= 32'hf979dc37;
8'h41 : rvCrc[11] <= 32'hfe8f3f31;
8'h42 : rvCrc[11] <= 32'hf6941a3b;
8'h43 : rvCrc[11] <= 32'hf162f93d;
8'h44 : rvCrc[11] <= 32'he6a2502f;
8'h45 : rvCrc[11] <= 32'he154b329;
8'h46 : rvCrc[11] <= 32'he94f9623;
8'h47 : rvCrc[11] <= 32'heeb97525;
8'h48 : rvCrc[11] <= 32'hc6cec407;
8'h49 : rvCrc[11] <= 32'hc1382701;
8'h4a : rvCrc[11] <= 32'hc923020b;
8'h4b : rvCrc[11] <= 32'hced5e10d;
8'h4c : rvCrc[11] <= 32'hd915481f;
8'h4d : rvCrc[11] <= 32'hdee3ab19;
8'h4e : rvCrc[11] <= 32'hd6f88e13;
8'h4f : rvCrc[11] <= 32'hd10e6d15;
8'h50 : rvCrc[11] <= 32'h8617ec57;
8'h51 : rvCrc[11] <= 32'h81e10f51;
8'h52 : rvCrc[11] <= 32'h89fa2a5b;
8'h53 : rvCrc[11] <= 32'h8e0cc95d;
8'h54 : rvCrc[11] <= 32'h99cc604f;
8'h55 : rvCrc[11] <= 32'h9e3a8349;
8'h56 : rvCrc[11] <= 32'h9621a643;
8'h57 : rvCrc[11] <= 32'h91d74545;
8'h58 : rvCrc[11] <= 32'hb9a0f467;
8'h59 : rvCrc[11] <= 32'hbe561761;
8'h5a : rvCrc[11] <= 32'hb64d326b;
8'h5b : rvCrc[11] <= 32'hb1bbd16d;
8'h5c : rvCrc[11] <= 32'ha67b787f;
8'h5d : rvCrc[11] <= 32'ha18d9b79;
8'h5e : rvCrc[11] <= 32'ha996be73;
8'h5f : rvCrc[11] <= 32'hae605d75;
8'h60 : rvCrc[11] <= 32'h07a5bcf7;
8'h61 : rvCrc[11] <= 32'h00535ff1;
8'h62 : rvCrc[11] <= 32'h08487afb;
8'h63 : rvCrc[11] <= 32'h0fbe99fd;
8'h64 : rvCrc[11] <= 32'h187e30ef;
8'h65 : rvCrc[11] <= 32'h1f88d3e9;
8'h66 : rvCrc[11] <= 32'h1793f6e3;
8'h67 : rvCrc[11] <= 32'h106515e5;
8'h68 : rvCrc[11] <= 32'h3812a4c7;
8'h69 : rvCrc[11] <= 32'h3fe447c1;
8'h6a : rvCrc[11] <= 32'h37ff62cb;
8'h6b : rvCrc[11] <= 32'h300981cd;
8'h6c : rvCrc[11] <= 32'h27c928df;
8'h6d : rvCrc[11] <= 32'h203fcbd9;
8'h6e : rvCrc[11] <= 32'h2824eed3;
8'h6f : rvCrc[11] <= 32'h2fd20dd5;
8'h70 : rvCrc[11] <= 32'h78cb8c97;
8'h71 : rvCrc[11] <= 32'h7f3d6f91;
8'h72 : rvCrc[11] <= 32'h77264a9b;
8'h73 : rvCrc[11] <= 32'h70d0a99d;
8'h74 : rvCrc[11] <= 32'h6710008f;
8'h75 : rvCrc[11] <= 32'h60e6e389;
8'h76 : rvCrc[11] <= 32'h68fdc683;
8'h77 : rvCrc[11] <= 32'h6f0b2585;
8'h78 : rvCrc[11] <= 32'h477c94a7;
8'h79 : rvCrc[11] <= 32'h408a77a1;
8'h7a : rvCrc[11] <= 32'h489152ab;
8'h7b : rvCrc[11] <= 32'h4f67b1ad;
8'h7c : rvCrc[11] <= 32'h58a718bf;
8'h7d : rvCrc[11] <= 32'h5f51fbb9;
8'h7e : rvCrc[11] <= 32'h574adeb3;
8'h7f : rvCrc[11] <= 32'h50bc3db5;
8'h80 : rvCrc[11] <= 32'hf632a5d9;
8'h81 : rvCrc[11] <= 32'hf1c446df;
8'h82 : rvCrc[11] <= 32'hf9df63d5;
8'h83 : rvCrc[11] <= 32'hfe2980d3;
8'h84 : rvCrc[11] <= 32'he9e929c1;
8'h85 : rvCrc[11] <= 32'hee1fcac7;
8'h86 : rvCrc[11] <= 32'he604efcd;
8'h87 : rvCrc[11] <= 32'he1f20ccb;
8'h88 : rvCrc[11] <= 32'hc985bde9;
8'h89 : rvCrc[11] <= 32'hce735eef;
8'h8a : rvCrc[11] <= 32'hc6687be5;
8'h8b : rvCrc[11] <= 32'hc19e98e3;
8'h8c : rvCrc[11] <= 32'hd65e31f1;
8'h8d : rvCrc[11] <= 32'hd1a8d2f7;
8'h8e : rvCrc[11] <= 32'hd9b3f7fd;
8'h8f : rvCrc[11] <= 32'hde4514fb;
8'h90 : rvCrc[11] <= 32'h895c95b9;
8'h91 : rvCrc[11] <= 32'h8eaa76bf;
8'h92 : rvCrc[11] <= 32'h86b153b5;
8'h93 : rvCrc[11] <= 32'h8147b0b3;
8'h94 : rvCrc[11] <= 32'h968719a1;
8'h95 : rvCrc[11] <= 32'h9171faa7;
8'h96 : rvCrc[11] <= 32'h996adfad;
8'h97 : rvCrc[11] <= 32'h9e9c3cab;
8'h98 : rvCrc[11] <= 32'hb6eb8d89;
8'h99 : rvCrc[11] <= 32'hb11d6e8f;
8'h9a : rvCrc[11] <= 32'hb9064b85;
8'h9b : rvCrc[11] <= 32'hbef0a883;
8'h9c : rvCrc[11] <= 32'ha9300191;
8'h9d : rvCrc[11] <= 32'haec6e297;
8'h9e : rvCrc[11] <= 32'ha6ddc79d;
8'h9f : rvCrc[11] <= 32'ha12b249b;
8'ha0 : rvCrc[11] <= 32'h08eec519;
8'ha1 : rvCrc[11] <= 32'h0f18261f;
8'ha2 : rvCrc[11] <= 32'h07030315;
8'ha3 : rvCrc[11] <= 32'h00f5e013;
8'ha4 : rvCrc[11] <= 32'h17354901;
8'ha5 : rvCrc[11] <= 32'h10c3aa07;
8'ha6 : rvCrc[11] <= 32'h18d88f0d;
8'ha7 : rvCrc[11] <= 32'h1f2e6c0b;
8'ha8 : rvCrc[11] <= 32'h3759dd29;
8'ha9 : rvCrc[11] <= 32'h30af3e2f;
8'haa : rvCrc[11] <= 32'h38b41b25;
8'hab : rvCrc[11] <= 32'h3f42f823;
8'hac : rvCrc[11] <= 32'h28825131;
8'had : rvCrc[11] <= 32'h2f74b237;
8'hae : rvCrc[11] <= 32'h276f973d;
8'haf : rvCrc[11] <= 32'h2099743b;
8'hb0 : rvCrc[11] <= 32'h7780f579;
8'hb1 : rvCrc[11] <= 32'h7076167f;
8'hb2 : rvCrc[11] <= 32'h786d3375;
8'hb3 : rvCrc[11] <= 32'h7f9bd073;
8'hb4 : rvCrc[11] <= 32'h685b7961;
8'hb5 : rvCrc[11] <= 32'h6fad9a67;
8'hb6 : rvCrc[11] <= 32'h67b6bf6d;
8'hb7 : rvCrc[11] <= 32'h60405c6b;
8'hb8 : rvCrc[11] <= 32'h4837ed49;
8'hb9 : rvCrc[11] <= 32'h4fc10e4f;
8'hba : rvCrc[11] <= 32'h47da2b45;
8'hbb : rvCrc[11] <= 32'h402cc843;
8'hbc : rvCrc[11] <= 32'h57ec6151;
8'hbd : rvCrc[11] <= 32'h501a8257;
8'hbe : rvCrc[11] <= 32'h5801a75d;
8'hbf : rvCrc[11] <= 32'h5ff7445b;
8'hc0 : rvCrc[11] <= 32'h0f4b79ee;
8'hc1 : rvCrc[11] <= 32'h08bd9ae8;
8'hc2 : rvCrc[11] <= 32'h00a6bfe2;
8'hc3 : rvCrc[11] <= 32'h07505ce4;
8'hc4 : rvCrc[11] <= 32'h1090f5f6;
8'hc5 : rvCrc[11] <= 32'h176616f0;
8'hc6 : rvCrc[11] <= 32'h1f7d33fa;
8'hc7 : rvCrc[11] <= 32'h188bd0fc;
8'hc8 : rvCrc[11] <= 32'h30fc61de;
8'hc9 : rvCrc[11] <= 32'h370a82d8;
8'hca : rvCrc[11] <= 32'h3f11a7d2;
8'hcb : rvCrc[11] <= 32'h38e744d4;
8'hcc : rvCrc[11] <= 32'h2f27edc6;
8'hcd : rvCrc[11] <= 32'h28d10ec0;
8'hce : rvCrc[11] <= 32'h20ca2bca;
8'hcf : rvCrc[11] <= 32'h273cc8cc;
8'hd0 : rvCrc[11] <= 32'h7025498e;
8'hd1 : rvCrc[11] <= 32'h77d3aa88;
8'hd2 : rvCrc[11] <= 32'h7fc88f82;
8'hd3 : rvCrc[11] <= 32'h783e6c84;
8'hd4 : rvCrc[11] <= 32'h6ffec596;
8'hd5 : rvCrc[11] <= 32'h68082690;
8'hd6 : rvCrc[11] <= 32'h6013039a;
8'hd7 : rvCrc[11] <= 32'h67e5e09c;
8'hd8 : rvCrc[11] <= 32'h4f9251be;
8'hd9 : rvCrc[11] <= 32'h4864b2b8;
8'hda : rvCrc[11] <= 32'h407f97b2;
8'hdb : rvCrc[11] <= 32'h478974b4;
8'hdc : rvCrc[11] <= 32'h5049dda6;
8'hdd : rvCrc[11] <= 32'h57bf3ea0;
8'hde : rvCrc[11] <= 32'h5fa41baa;
8'hdf : rvCrc[11] <= 32'h5852f8ac;
8'he0 : rvCrc[11] <= 32'hf197192e;
8'he1 : rvCrc[11] <= 32'hf661fa28;
8'he2 : rvCrc[11] <= 32'hfe7adf22;
8'he3 : rvCrc[11] <= 32'hf98c3c24;
8'he4 : rvCrc[11] <= 32'hee4c9536;
8'he5 : rvCrc[11] <= 32'he9ba7630;
8'he6 : rvCrc[11] <= 32'he1a1533a;
8'he7 : rvCrc[11] <= 32'he657b03c;
8'he8 : rvCrc[11] <= 32'hce20011e;
8'he9 : rvCrc[11] <= 32'hc9d6e218;
8'hea : rvCrc[11] <= 32'hc1cdc712;
8'heb : rvCrc[11] <= 32'hc63b2414;
8'hec : rvCrc[11] <= 32'hd1fb8d06;
8'hed : rvCrc[11] <= 32'hd60d6e00;
8'hee : rvCrc[11] <= 32'hde164b0a;
8'hef : rvCrc[11] <= 32'hd9e0a80c;
8'hf0 : rvCrc[11] <= 32'h8ef9294e;
8'hf1 : rvCrc[11] <= 32'h890fca48;
8'hf2 : rvCrc[11] <= 32'h8114ef42;
8'hf3 : rvCrc[11] <= 32'h86e20c44;
8'hf4 : rvCrc[11] <= 32'h9122a556;
8'hf5 : rvCrc[11] <= 32'h96d44650;
8'hf6 : rvCrc[11] <= 32'h9ecf635a;
8'hf7 : rvCrc[11] <= 32'h9939805c;
8'hf8 : rvCrc[11] <= 32'hb14e317e;
8'hf9 : rvCrc[11] <= 32'hb6b8d278;
8'hfa : rvCrc[11] <= 32'hbea3f772;
8'hfb : rvCrc[11] <= 32'hb9551474;
8'hfc : rvCrc[11] <= 32'hae95bd66;
8'hfd : rvCrc[11] <= 32'ha9635e60;
8'hfe : rvCrc[11] <= 32'ha1787b6a;
8'hff : rvCrc[11] <= 32'ha68e986c;
endcase
case(iv_Input[103:096])
8'h00 : rvCrc[12] <= 32'h00000000;
8'h01 : rvCrc[12] <= 32'he8a45605;
8'h02 : rvCrc[12] <= 32'hd589b1bd;
8'h03 : rvCrc[12] <= 32'h3d2de7b8;
8'h04 : rvCrc[12] <= 32'hafd27ecd;
8'h05 : rvCrc[12] <= 32'h477628c8;
8'h06 : rvCrc[12] <= 32'h7a5bcf70;
8'h07 : rvCrc[12] <= 32'h92ff9975;
8'h08 : rvCrc[12] <= 32'h5b65e02d;
8'h09 : rvCrc[12] <= 32'hb3c1b628;
8'h0a : rvCrc[12] <= 32'h8eec5190;
8'h0b : rvCrc[12] <= 32'h66480795;
8'h0c : rvCrc[12] <= 32'hf4b79ee0;
8'h0d : rvCrc[12] <= 32'h1c13c8e5;
8'h0e : rvCrc[12] <= 32'h213e2f5d;
8'h0f : rvCrc[12] <= 32'hc99a7958;
8'h10 : rvCrc[12] <= 32'hb6cbc05a;
8'h11 : rvCrc[12] <= 32'h5e6f965f;
8'h12 : rvCrc[12] <= 32'h634271e7;
8'h13 : rvCrc[12] <= 32'h8be627e2;
8'h14 : rvCrc[12] <= 32'h1919be97;
8'h15 : rvCrc[12] <= 32'hf1bde892;
8'h16 : rvCrc[12] <= 32'hcc900f2a;
8'h17 : rvCrc[12] <= 32'h2434592f;
8'h18 : rvCrc[12] <= 32'hedae2077;
8'h19 : rvCrc[12] <= 32'h050a7672;
8'h1a : rvCrc[12] <= 32'h382791ca;
8'h1b : rvCrc[12] <= 32'hd083c7cf;
8'h1c : rvCrc[12] <= 32'h427c5eba;
8'h1d : rvCrc[12] <= 32'haad808bf;
8'h1e : rvCrc[12] <= 32'h97f5ef07;
8'h1f : rvCrc[12] <= 32'h7f51b902;
8'h20 : rvCrc[12] <= 32'h69569d03;
8'h21 : rvCrc[12] <= 32'h81f2cb06;
8'h22 : rvCrc[12] <= 32'hbcdf2cbe;
8'h23 : rvCrc[12] <= 32'h547b7abb;
8'h24 : rvCrc[12] <= 32'hc684e3ce;
8'h25 : rvCrc[12] <= 32'h2e20b5cb;
8'h26 : rvCrc[12] <= 32'h130d5273;
8'h27 : rvCrc[12] <= 32'hfba90476;
8'h28 : rvCrc[12] <= 32'h32337d2e;
8'h29 : rvCrc[12] <= 32'hda972b2b;
8'h2a : rvCrc[12] <= 32'he7bacc93;
8'h2b : rvCrc[12] <= 32'h0f1e9a96;
8'h2c : rvCrc[12] <= 32'h9de103e3;
8'h2d : rvCrc[12] <= 32'h754555e6;
8'h2e : rvCrc[12] <= 32'h4868b25e;
8'h2f : rvCrc[12] <= 32'ha0cce45b;
8'h30 : rvCrc[12] <= 32'hdf9d5d59;
8'h31 : rvCrc[12] <= 32'h37390b5c;
8'h32 : rvCrc[12] <= 32'h0a14ece4;
8'h33 : rvCrc[12] <= 32'he2b0bae1;
8'h34 : rvCrc[12] <= 32'h704f2394;
8'h35 : rvCrc[12] <= 32'h98eb7591;
8'h36 : rvCrc[12] <= 32'ha5c69229;
8'h37 : rvCrc[12] <= 32'h4d62c42c;
8'h38 : rvCrc[12] <= 32'h84f8bd74;
8'h39 : rvCrc[12] <= 32'h6c5ceb71;
8'h3a : rvCrc[12] <= 32'h51710cc9;
8'h3b : rvCrc[12] <= 32'hb9d55acc;
8'h3c : rvCrc[12] <= 32'h2b2ac3b9;
8'h3d : rvCrc[12] <= 32'hc38e95bc;
8'h3e : rvCrc[12] <= 32'hfea37204;
8'h3f : rvCrc[12] <= 32'h16072401;
8'h40 : rvCrc[12] <= 32'hd2ad3a06;
8'h41 : rvCrc[12] <= 32'h3a096c03;
8'h42 : rvCrc[12] <= 32'h07248bbb;
8'h43 : rvCrc[12] <= 32'hef80ddbe;
8'h44 : rvCrc[12] <= 32'h7d7f44cb;
8'h45 : rvCrc[12] <= 32'h95db12ce;
8'h46 : rvCrc[12] <= 32'ha8f6f576;
8'h47 : rvCrc[12] <= 32'h4052a373;
8'h48 : rvCrc[12] <= 32'h89c8da2b;
8'h49 : rvCrc[12] <= 32'h616c8c2e;
8'h4a : rvCrc[12] <= 32'h5c416b96;
8'h4b : rvCrc[12] <= 32'hb4e53d93;
8'h4c : rvCrc[12] <= 32'h261aa4e6;
8'h4d : rvCrc[12] <= 32'hcebef2e3;
8'h4e : rvCrc[12] <= 32'hf393155b;
8'h4f : rvCrc[12] <= 32'h1b37435e;
8'h50 : rvCrc[12] <= 32'h6466fa5c;
8'h51 : rvCrc[12] <= 32'h8cc2ac59;
8'h52 : rvCrc[12] <= 32'hb1ef4be1;
8'h53 : rvCrc[12] <= 32'h594b1de4;
8'h54 : rvCrc[12] <= 32'hcbb48491;
8'h55 : rvCrc[12] <= 32'h2310d294;
8'h56 : rvCrc[12] <= 32'h1e3d352c;
8'h57 : rvCrc[12] <= 32'hf6996329;
8'h58 : rvCrc[12] <= 32'h3f031a71;
8'h59 : rvCrc[12] <= 32'hd7a74c74;
8'h5a : rvCrc[12] <= 32'hea8aabcc;
8'h5b : rvCrc[12] <= 32'h022efdc9;
8'h5c : rvCrc[12] <= 32'h90d164bc;
8'h5d : rvCrc[12] <= 32'h787532b9;
8'h5e : rvCrc[12] <= 32'h4558d501;
8'h5f : rvCrc[12] <= 32'hadfc8304;
8'h60 : rvCrc[12] <= 32'hbbfba705;
8'h61 : rvCrc[12] <= 32'h535ff100;
8'h62 : rvCrc[12] <= 32'h6e7216b8;
8'h63 : rvCrc[12] <= 32'h86d640bd;
8'h64 : rvCrc[12] <= 32'h1429d9c8;
8'h65 : rvCrc[12] <= 32'hfc8d8fcd;
8'h66 : rvCrc[12] <= 32'hc1a06875;
8'h67 : rvCrc[12] <= 32'h29043e70;
8'h68 : rvCrc[12] <= 32'he09e4728;
8'h69 : rvCrc[12] <= 32'h083a112d;
8'h6a : rvCrc[12] <= 32'h3517f695;
8'h6b : rvCrc[12] <= 32'hddb3a090;
8'h6c : rvCrc[12] <= 32'h4f4c39e5;
8'h6d : rvCrc[12] <= 32'ha7e86fe0;
8'h6e : rvCrc[12] <= 32'h9ac58858;
8'h6f : rvCrc[12] <= 32'h7261de5d;
8'h70 : rvCrc[12] <= 32'h0d30675f;
8'h71 : rvCrc[12] <= 32'he594315a;
8'h72 : rvCrc[12] <= 32'hd8b9d6e2;
8'h73 : rvCrc[12] <= 32'h301d80e7;
8'h74 : rvCrc[12] <= 32'ha2e21992;
8'h75 : rvCrc[12] <= 32'h4a464f97;
8'h76 : rvCrc[12] <= 32'h776ba82f;
8'h77 : rvCrc[12] <= 32'h9fcffe2a;
8'h78 : rvCrc[12] <= 32'h56558772;
8'h79 : rvCrc[12] <= 32'hbef1d177;
8'h7a : rvCrc[12] <= 32'h83dc36cf;
8'h7b : rvCrc[12] <= 32'h6b7860ca;
8'h7c : rvCrc[12] <= 32'hf987f9bf;
8'h7d : rvCrc[12] <= 32'h1123afba;
8'h7e : rvCrc[12] <= 32'h2c0e4802;
8'h7f : rvCrc[12] <= 32'hc4aa1e07;
8'h80 : rvCrc[12] <= 32'ha19b69bb;
8'h81 : rvCrc[12] <= 32'h493f3fbe;
8'h82 : rvCrc[12] <= 32'h7412d806;
8'h83 : rvCrc[12] <= 32'h9cb68e03;
8'h84 : rvCrc[12] <= 32'h0e491776;
8'h85 : rvCrc[12] <= 32'he6ed4173;
8'h86 : rvCrc[12] <= 32'hdbc0a6cb;
8'h87 : rvCrc[12] <= 32'h3364f0ce;
8'h88 : rvCrc[12] <= 32'hfafe8996;
8'h89 : rvCrc[12] <= 32'h125adf93;
8'h8a : rvCrc[12] <= 32'h2f77382b;
8'h8b : rvCrc[12] <= 32'hc7d36e2e;
8'h8c : rvCrc[12] <= 32'h552cf75b;
8'h8d : rvCrc[12] <= 32'hbd88a15e;
8'h8e : rvCrc[12] <= 32'h80a546e6;
8'h8f : rvCrc[12] <= 32'h680110e3;
8'h90 : rvCrc[12] <= 32'h1750a9e1;
8'h91 : rvCrc[12] <= 32'hfff4ffe4;
8'h92 : rvCrc[12] <= 32'hc2d9185c;
8'h93 : rvCrc[12] <= 32'h2a7d4e59;
8'h94 : rvCrc[12] <= 32'hb882d72c;
8'h95 : rvCrc[12] <= 32'h50268129;
8'h96 : rvCrc[12] <= 32'h6d0b6691;
8'h97 : rvCrc[12] <= 32'h85af3094;
8'h98 : rvCrc[12] <= 32'h4c3549cc;
8'h99 : rvCrc[12] <= 32'ha4911fc9;
8'h9a : rvCrc[12] <= 32'h99bcf871;
8'h9b : rvCrc[12] <= 32'h7118ae74;
8'h9c : rvCrc[12] <= 32'he3e73701;
8'h9d : rvCrc[12] <= 32'h0b436104;
8'h9e : rvCrc[12] <= 32'h366e86bc;
8'h9f : rvCrc[12] <= 32'hdecad0b9;
8'ha0 : rvCrc[12] <= 32'hc8cdf4b8;
8'ha1 : rvCrc[12] <= 32'h2069a2bd;
8'ha2 : rvCrc[12] <= 32'h1d444505;
8'ha3 : rvCrc[12] <= 32'hf5e01300;
8'ha4 : rvCrc[12] <= 32'h671f8a75;
8'ha5 : rvCrc[12] <= 32'h8fbbdc70;
8'ha6 : rvCrc[12] <= 32'hb2963bc8;
8'ha7 : rvCrc[12] <= 32'h5a326dcd;
8'ha8 : rvCrc[12] <= 32'h93a81495;
8'ha9 : rvCrc[12] <= 32'h7b0c4290;
8'haa : rvCrc[12] <= 32'h4621a528;
8'hab : rvCrc[12] <= 32'hae85f32d;
8'hac : rvCrc[12] <= 32'h3c7a6a58;
8'had : rvCrc[12] <= 32'hd4de3c5d;
8'hae : rvCrc[12] <= 32'he9f3dbe5;
8'haf : rvCrc[12] <= 32'h01578de0;
8'hb0 : rvCrc[12] <= 32'h7e0634e2;
8'hb1 : rvCrc[12] <= 32'h96a262e7;
8'hb2 : rvCrc[12] <= 32'hab8f855f;
8'hb3 : rvCrc[12] <= 32'h432bd35a;
8'hb4 : rvCrc[12] <= 32'hd1d44a2f;
8'hb5 : rvCrc[12] <= 32'h39701c2a;
8'hb6 : rvCrc[12] <= 32'h045dfb92;
8'hb7 : rvCrc[12] <= 32'hecf9ad97;
8'hb8 : rvCrc[12] <= 32'h2563d4cf;
8'hb9 : rvCrc[12] <= 32'hcdc782ca;
8'hba : rvCrc[12] <= 32'hf0ea6572;
8'hbb : rvCrc[12] <= 32'h184e3377;
8'hbc : rvCrc[12] <= 32'h8ab1aa02;
8'hbd : rvCrc[12] <= 32'h6215fc07;
8'hbe : rvCrc[12] <= 32'h5f381bbf;
8'hbf : rvCrc[12] <= 32'hb79c4dba;
8'hc0 : rvCrc[12] <= 32'h733653bd;
8'hc1 : rvCrc[12] <= 32'h9b9205b8;
8'hc2 : rvCrc[12] <= 32'ha6bfe200;
8'hc3 : rvCrc[12] <= 32'h4e1bb405;
8'hc4 : rvCrc[12] <= 32'hdce42d70;
8'hc5 : rvCrc[12] <= 32'h34407b75;
8'hc6 : rvCrc[12] <= 32'h096d9ccd;
8'hc7 : rvCrc[12] <= 32'he1c9cac8;
8'hc8 : rvCrc[12] <= 32'h2853b390;
8'hc9 : rvCrc[12] <= 32'hc0f7e595;
8'hca : rvCrc[12] <= 32'hfdda022d;
8'hcb : rvCrc[12] <= 32'h157e5428;
8'hcc : rvCrc[12] <= 32'h8781cd5d;
8'hcd : rvCrc[12] <= 32'h6f259b58;
8'hce : rvCrc[12] <= 32'h52087ce0;
8'hcf : rvCrc[12] <= 32'hbaac2ae5;
8'hd0 : rvCrc[12] <= 32'hc5fd93e7;
8'hd1 : rvCrc[12] <= 32'h2d59c5e2;
8'hd2 : rvCrc[12] <= 32'h1074225a;
8'hd3 : rvCrc[12] <= 32'hf8d0745f;
8'hd4 : rvCrc[12] <= 32'h6a2fed2a;
8'hd5 : rvCrc[12] <= 32'h828bbb2f;
8'hd6 : rvCrc[12] <= 32'hbfa65c97;
8'hd7 : rvCrc[12] <= 32'h57020a92;
8'hd8 : rvCrc[12] <= 32'h9e9873ca;
8'hd9 : rvCrc[12] <= 32'h763c25cf;
8'hda : rvCrc[12] <= 32'h4b11c277;
8'hdb : rvCrc[12] <= 32'ha3b59472;
8'hdc : rvCrc[12] <= 32'h314a0d07;
8'hdd : rvCrc[12] <= 32'hd9ee5b02;
8'hde : rvCrc[12] <= 32'he4c3bcba;
8'hdf : rvCrc[12] <= 32'h0c67eabf;
8'he0 : rvCrc[12] <= 32'h1a60cebe;
8'he1 : rvCrc[12] <= 32'hf2c498bb;
8'he2 : rvCrc[12] <= 32'hcfe97f03;
8'he3 : rvCrc[12] <= 32'h274d2906;
8'he4 : rvCrc[12] <= 32'hb5b2b073;
8'he5 : rvCrc[12] <= 32'h5d16e676;
8'he6 : rvCrc[12] <= 32'h603b01ce;
8'he7 : rvCrc[12] <= 32'h889f57cb;
8'he8 : rvCrc[12] <= 32'h41052e93;
8'he9 : rvCrc[12] <= 32'ha9a17896;
8'hea : rvCrc[12] <= 32'h948c9f2e;
8'heb : rvCrc[12] <= 32'h7c28c92b;
8'hec : rvCrc[12] <= 32'heed7505e;
8'hed : rvCrc[12] <= 32'h0673065b;
8'hee : rvCrc[12] <= 32'h3b5ee1e3;
8'hef : rvCrc[12] <= 32'hd3fab7e6;
8'hf0 : rvCrc[12] <= 32'hacab0ee4;
8'hf1 : rvCrc[12] <= 32'h440f58e1;
8'hf2 : rvCrc[12] <= 32'h7922bf59;
8'hf3 : rvCrc[12] <= 32'h9186e95c;
8'hf4 : rvCrc[12] <= 32'h03797029;
8'hf5 : rvCrc[12] <= 32'hebdd262c;
8'hf6 : rvCrc[12] <= 32'hd6f0c194;
8'hf7 : rvCrc[12] <= 32'h3e549791;
8'hf8 : rvCrc[12] <= 32'hf7ceeec9;
8'hf9 : rvCrc[12] <= 32'h1f6ab8cc;
8'hfa : rvCrc[12] <= 32'h22475f74;
8'hfb : rvCrc[12] <= 32'hcae30971;
8'hfc : rvCrc[12] <= 32'h581c9004;
8'hfd : rvCrc[12] <= 32'hb0b8c601;
8'hfe : rvCrc[12] <= 32'h8d9521b9;
8'hff : rvCrc[12] <= 32'h653177bc;
endcase
case(iv_Input[111:104])
8'h00 : rvCrc[13] <= 32'h00000000;
8'h01 : rvCrc[13] <= 32'h47f7cec1;
8'h02 : rvCrc[13] <= 32'h8fef9d82;
8'h03 : rvCrc[13] <= 32'hc8185343;
8'h04 : rvCrc[13] <= 32'h1b1e26b3;
8'h05 : rvCrc[13] <= 32'h5ce9e872;
8'h06 : rvCrc[13] <= 32'h94f1bb31;
8'h07 : rvCrc[13] <= 32'hd30675f0;
8'h08 : rvCrc[13] <= 32'h363c4d66;
8'h09 : rvCrc[13] <= 32'h71cb83a7;
8'h0a : rvCrc[13] <= 32'hb9d3d0e4;
8'h0b : rvCrc[13] <= 32'hfe241e25;
8'h0c : rvCrc[13] <= 32'h2d226bd5;
8'h0d : rvCrc[13] <= 32'h6ad5a514;
8'h0e : rvCrc[13] <= 32'ha2cdf657;
8'h0f : rvCrc[13] <= 32'he53a3896;
8'h10 : rvCrc[13] <= 32'h6c789acc;
8'h11 : rvCrc[13] <= 32'h2b8f540d;
8'h12 : rvCrc[13] <= 32'he397074e;
8'h13 : rvCrc[13] <= 32'ha460c98f;
8'h14 : rvCrc[13] <= 32'h7766bc7f;
8'h15 : rvCrc[13] <= 32'h309172be;
8'h16 : rvCrc[13] <= 32'hf88921fd;
8'h17 : rvCrc[13] <= 32'hbf7eef3c;
8'h18 : rvCrc[13] <= 32'h5a44d7aa;
8'h19 : rvCrc[13] <= 32'h1db3196b;
8'h1a : rvCrc[13] <= 32'hd5ab4a28;
8'h1b : rvCrc[13] <= 32'h925c84e9;
8'h1c : rvCrc[13] <= 32'h415af119;
8'h1d : rvCrc[13] <= 32'h06ad3fd8;
8'h1e : rvCrc[13] <= 32'hceb56c9b;
8'h1f : rvCrc[13] <= 32'h8942a25a;
8'h20 : rvCrc[13] <= 32'hd8f13598;
8'h21 : rvCrc[13] <= 32'h9f06fb59;
8'h22 : rvCrc[13] <= 32'h571ea81a;
8'h23 : rvCrc[13] <= 32'h10e966db;
8'h24 : rvCrc[13] <= 32'hc3ef132b;
8'h25 : rvCrc[13] <= 32'h8418ddea;
8'h26 : rvCrc[13] <= 32'h4c008ea9;
8'h27 : rvCrc[13] <= 32'h0bf74068;
8'h28 : rvCrc[13] <= 32'heecd78fe;
8'h29 : rvCrc[13] <= 32'ha93ab63f;
8'h2a : rvCrc[13] <= 32'h6122e57c;
8'h2b : rvCrc[13] <= 32'h26d52bbd;
8'h2c : rvCrc[13] <= 32'hf5d35e4d;
8'h2d : rvCrc[13] <= 32'hb224908c;
8'h2e : rvCrc[13] <= 32'h7a3cc3cf;
8'h2f : rvCrc[13] <= 32'h3dcb0d0e;
8'h30 : rvCrc[13] <= 32'hb489af54;
8'h31 : rvCrc[13] <= 32'hf37e6195;
8'h32 : rvCrc[13] <= 32'h3b6632d6;
8'h33 : rvCrc[13] <= 32'h7c91fc17;
8'h34 : rvCrc[13] <= 32'haf9789e7;
8'h35 : rvCrc[13] <= 32'he8604726;
8'h36 : rvCrc[13] <= 32'h20781465;
8'h37 : rvCrc[13] <= 32'h678fdaa4;
8'h38 : rvCrc[13] <= 32'h82b5e232;
8'h39 : rvCrc[13] <= 32'hc5422cf3;
8'h3a : rvCrc[13] <= 32'h0d5a7fb0;
8'h3b : rvCrc[13] <= 32'h4aadb171;
8'h3c : rvCrc[13] <= 32'h99abc481;
8'h3d : rvCrc[13] <= 32'hde5c0a40;
8'h3e : rvCrc[13] <= 32'h16445903;
8'h3f : rvCrc[13] <= 32'h51b397c2;
8'h40 : rvCrc[13] <= 32'hb5237687;
8'h41 : rvCrc[13] <= 32'hf2d4b846;
8'h42 : rvCrc[13] <= 32'h3acceb05;
8'h43 : rvCrc[13] <= 32'h7d3b25c4;
8'h44 : rvCrc[13] <= 32'hae3d5034;
8'h45 : rvCrc[13] <= 32'he9ca9ef5;
8'h46 : rvCrc[13] <= 32'h21d2cdb6;
8'h47 : rvCrc[13] <= 32'h66250377;
8'h48 : rvCrc[13] <= 32'h831f3be1;
8'h49 : rvCrc[13] <= 32'hc4e8f520;
8'h4a : rvCrc[13] <= 32'h0cf0a663;
8'h4b : rvCrc[13] <= 32'h4b0768a2;
8'h4c : rvCrc[13] <= 32'h98011d52;
8'h4d : rvCrc[13] <= 32'hdff6d393;
8'h4e : rvCrc[13] <= 32'h17ee80d0;
8'h4f : rvCrc[13] <= 32'h50194e11;
8'h50 : rvCrc[13] <= 32'hd95bec4b;
8'h51 : rvCrc[13] <= 32'h9eac228a;
8'h52 : rvCrc[13] <= 32'h56b471c9;
8'h53 : rvCrc[13] <= 32'h1143bf08;
8'h54 : rvCrc[13] <= 32'hc245caf8;
8'h55 : rvCrc[13] <= 32'h85b20439;
8'h56 : rvCrc[13] <= 32'h4daa577a;
8'h57 : rvCrc[13] <= 32'h0a5d99bb;
8'h58 : rvCrc[13] <= 32'hef67a12d;
8'h59 : rvCrc[13] <= 32'ha8906fec;
8'h5a : rvCrc[13] <= 32'h60883caf;
8'h5b : rvCrc[13] <= 32'h277ff26e;
8'h5c : rvCrc[13] <= 32'hf479879e;
8'h5d : rvCrc[13] <= 32'hb38e495f;
8'h5e : rvCrc[13] <= 32'h7b961a1c;
8'h5f : rvCrc[13] <= 32'h3c61d4dd;
8'h60 : rvCrc[13] <= 32'h6dd2431f;
8'h61 : rvCrc[13] <= 32'h2a258dde;
8'h62 : rvCrc[13] <= 32'he23dde9d;
8'h63 : rvCrc[13] <= 32'ha5ca105c;
8'h64 : rvCrc[13] <= 32'h76cc65ac;
8'h65 : rvCrc[13] <= 32'h313bab6d;
8'h66 : rvCrc[13] <= 32'hf923f82e;
8'h67 : rvCrc[13] <= 32'hbed436ef;
8'h68 : rvCrc[13] <= 32'h5bee0e79;
8'h69 : rvCrc[13] <= 32'h1c19c0b8;
8'h6a : rvCrc[13] <= 32'hd40193fb;
8'h6b : rvCrc[13] <= 32'h93f65d3a;
8'h6c : rvCrc[13] <= 32'h40f028ca;
8'h6d : rvCrc[13] <= 32'h0707e60b;
8'h6e : rvCrc[13] <= 32'hcf1fb548;
8'h6f : rvCrc[13] <= 32'h88e87b89;
8'h70 : rvCrc[13] <= 32'h01aad9d3;
8'h71 : rvCrc[13] <= 32'h465d1712;
8'h72 : rvCrc[13] <= 32'h8e454451;
8'h73 : rvCrc[13] <= 32'hc9b28a90;
8'h74 : rvCrc[13] <= 32'h1ab4ff60;
8'h75 : rvCrc[13] <= 32'h5d4331a1;
8'h76 : rvCrc[13] <= 32'h955b62e2;
8'h77 : rvCrc[13] <= 32'hd2acac23;
8'h78 : rvCrc[13] <= 32'h379694b5;
8'h79 : rvCrc[13] <= 32'h70615a74;
8'h7a : rvCrc[13] <= 32'hb8790937;
8'h7b : rvCrc[13] <= 32'hff8ec7f6;
8'h7c : rvCrc[13] <= 32'h2c88b206;
8'h7d : rvCrc[13] <= 32'h6b7f7cc7;
8'h7e : rvCrc[13] <= 32'ha3672f84;
8'h7f : rvCrc[13] <= 32'he490e145;
8'h80 : rvCrc[13] <= 32'h6e87f0b9;
8'h81 : rvCrc[13] <= 32'h29703e78;
8'h82 : rvCrc[13] <= 32'he1686d3b;
8'h83 : rvCrc[13] <= 32'ha69fa3fa;
8'h84 : rvCrc[13] <= 32'h7599d60a;
8'h85 : rvCrc[13] <= 32'h326e18cb;
8'h86 : rvCrc[13] <= 32'hfa764b88;
8'h87 : rvCrc[13] <= 32'hbd818549;
8'h88 : rvCrc[13] <= 32'h58bbbddf;
8'h89 : rvCrc[13] <= 32'h1f4c731e;
8'h8a : rvCrc[13] <= 32'hd754205d;
8'h8b : rvCrc[13] <= 32'h90a3ee9c;
8'h8c : rvCrc[13] <= 32'h43a59b6c;
8'h8d : rvCrc[13] <= 32'h045255ad;
8'h8e : rvCrc[13] <= 32'hcc4a06ee;
8'h8f : rvCrc[13] <= 32'h8bbdc82f;
8'h90 : rvCrc[13] <= 32'h02ff6a75;
8'h91 : rvCrc[13] <= 32'h4508a4b4;
8'h92 : rvCrc[13] <= 32'h8d10f7f7;
8'h93 : rvCrc[13] <= 32'hcae73936;
8'h94 : rvCrc[13] <= 32'h19e14cc6;
8'h95 : rvCrc[13] <= 32'h5e168207;
8'h96 : rvCrc[13] <= 32'h960ed144;
8'h97 : rvCrc[13] <= 32'hd1f91f85;
8'h98 : rvCrc[13] <= 32'h34c32713;
8'h99 : rvCrc[13] <= 32'h7334e9d2;
8'h9a : rvCrc[13] <= 32'hbb2cba91;
8'h9b : rvCrc[13] <= 32'hfcdb7450;
8'h9c : rvCrc[13] <= 32'h2fdd01a0;
8'h9d : rvCrc[13] <= 32'h682acf61;
8'h9e : rvCrc[13] <= 32'ha0329c22;
8'h9f : rvCrc[13] <= 32'he7c552e3;
8'ha0 : rvCrc[13] <= 32'hb676c521;
8'ha1 : rvCrc[13] <= 32'hf1810be0;
8'ha2 : rvCrc[13] <= 32'h399958a3;
8'ha3 : rvCrc[13] <= 32'h7e6e9662;
8'ha4 : rvCrc[13] <= 32'had68e392;
8'ha5 : rvCrc[13] <= 32'hea9f2d53;
8'ha6 : rvCrc[13] <= 32'h22877e10;
8'ha7 : rvCrc[13] <= 32'h6570b0d1;
8'ha8 : rvCrc[13] <= 32'h804a8847;
8'ha9 : rvCrc[13] <= 32'hc7bd4686;
8'haa : rvCrc[13] <= 32'h0fa515c5;
8'hab : rvCrc[13] <= 32'h4852db04;
8'hac : rvCrc[13] <= 32'h9b54aef4;
8'had : rvCrc[13] <= 32'hdca36035;
8'hae : rvCrc[13] <= 32'h14bb3376;
8'haf : rvCrc[13] <= 32'h534cfdb7;
8'hb0 : rvCrc[13] <= 32'hda0e5fed;
8'hb1 : rvCrc[13] <= 32'h9df9912c;
8'hb2 : rvCrc[13] <= 32'h55e1c26f;
8'hb3 : rvCrc[13] <= 32'h12160cae;
8'hb4 : rvCrc[13] <= 32'hc110795e;
8'hb5 : rvCrc[13] <= 32'h86e7b79f;
8'hb6 : rvCrc[13] <= 32'h4effe4dc;
8'hb7 : rvCrc[13] <= 32'h09082a1d;
8'hb8 : rvCrc[13] <= 32'hec32128b;
8'hb9 : rvCrc[13] <= 32'habc5dc4a;
8'hba : rvCrc[13] <= 32'h63dd8f09;
8'hbb : rvCrc[13] <= 32'h242a41c8;
8'hbc : rvCrc[13] <= 32'hf72c3438;
8'hbd : rvCrc[13] <= 32'hb0dbfaf9;
8'hbe : rvCrc[13] <= 32'h78c3a9ba;
8'hbf : rvCrc[13] <= 32'h3f34677b;
8'hc0 : rvCrc[13] <= 32'hdba4863e;
8'hc1 : rvCrc[13] <= 32'h9c5348ff;
8'hc2 : rvCrc[13] <= 32'h544b1bbc;
8'hc3 : rvCrc[13] <= 32'h13bcd57d;
8'hc4 : rvCrc[13] <= 32'hc0baa08d;
8'hc5 : rvCrc[13] <= 32'h874d6e4c;
8'hc6 : rvCrc[13] <= 32'h4f553d0f;
8'hc7 : rvCrc[13] <= 32'h08a2f3ce;
8'hc8 : rvCrc[13] <= 32'hed98cb58;
8'hc9 : rvCrc[13] <= 32'haa6f0599;
8'hca : rvCrc[13] <= 32'h627756da;
8'hcb : rvCrc[13] <= 32'h2580981b;
8'hcc : rvCrc[13] <= 32'hf686edeb;
8'hcd : rvCrc[13] <= 32'hb171232a;
8'hce : rvCrc[13] <= 32'h79697069;
8'hcf : rvCrc[13] <= 32'h3e9ebea8;
8'hd0 : rvCrc[13] <= 32'hb7dc1cf2;
8'hd1 : rvCrc[13] <= 32'hf02bd233;
8'hd2 : rvCrc[13] <= 32'h38338170;
8'hd3 : rvCrc[13] <= 32'h7fc44fb1;
8'hd4 : rvCrc[13] <= 32'hacc23a41;
8'hd5 : rvCrc[13] <= 32'heb35f480;
8'hd6 : rvCrc[13] <= 32'h232da7c3;
8'hd7 : rvCrc[13] <= 32'h64da6902;
8'hd8 : rvCrc[13] <= 32'h81e05194;
8'hd9 : rvCrc[13] <= 32'hc6179f55;
8'hda : rvCrc[13] <= 32'h0e0fcc16;
8'hdb : rvCrc[13] <= 32'h49f802d7;
8'hdc : rvCrc[13] <= 32'h9afe7727;
8'hdd : rvCrc[13] <= 32'hdd09b9e6;
8'hde : rvCrc[13] <= 32'h1511eaa5;
8'hdf : rvCrc[13] <= 32'h52e62464;
8'he0 : rvCrc[13] <= 32'h0355b3a6;
8'he1 : rvCrc[13] <= 32'h44a27d67;
8'he2 : rvCrc[13] <= 32'h8cba2e24;
8'he3 : rvCrc[13] <= 32'hcb4de0e5;
8'he4 : rvCrc[13] <= 32'h184b9515;
8'he5 : rvCrc[13] <= 32'h5fbc5bd4;
8'he6 : rvCrc[13] <= 32'h97a40897;
8'he7 : rvCrc[13] <= 32'hd053c656;
8'he8 : rvCrc[13] <= 32'h3569fec0;
8'he9 : rvCrc[13] <= 32'h729e3001;
8'hea : rvCrc[13] <= 32'hba866342;
8'heb : rvCrc[13] <= 32'hfd71ad83;
8'hec : rvCrc[13] <= 32'h2e77d873;
8'hed : rvCrc[13] <= 32'h698016b2;
8'hee : rvCrc[13] <= 32'ha19845f1;
8'hef : rvCrc[13] <= 32'he66f8b30;
8'hf0 : rvCrc[13] <= 32'h6f2d296a;
8'hf1 : rvCrc[13] <= 32'h28dae7ab;
8'hf2 : rvCrc[13] <= 32'he0c2b4e8;
8'hf3 : rvCrc[13] <= 32'ha7357a29;
8'hf4 : rvCrc[13] <= 32'h74330fd9;
8'hf5 : rvCrc[13] <= 32'h33c4c118;
8'hf6 : rvCrc[13] <= 32'hfbdc925b;
8'hf7 : rvCrc[13] <= 32'hbc2b5c9a;
8'hf8 : rvCrc[13] <= 32'h5911640c;
8'hf9 : rvCrc[13] <= 32'h1ee6aacd;
8'hfa : rvCrc[13] <= 32'hd6fef98e;
8'hfb : rvCrc[13] <= 32'h9109374f;
8'hfc : rvCrc[13] <= 32'h420f42bf;
8'hfd : rvCrc[13] <= 32'h05f88c7e;
8'hfe : rvCrc[13] <= 32'hcde0df3d;
8'hff : rvCrc[13] <= 32'h8a1711fc;
endcase
case(iv_Input[119:112])
8'h00 : rvCrc[14] <= 32'h00000000;
8'h01 : rvCrc[14] <= 32'hdd0fe172;
8'h02 : rvCrc[14] <= 32'hbededf53;
8'h03 : rvCrc[14] <= 32'h63d13e21;
8'h04 : rvCrc[14] <= 32'h797ca311;
8'h05 : rvCrc[14] <= 32'ha4734263;
8'h06 : rvCrc[14] <= 32'hc7a27c42;
8'h07 : rvCrc[14] <= 32'h1aad9d30;
8'h08 : rvCrc[14] <= 32'hf2f94622;
8'h09 : rvCrc[14] <= 32'h2ff6a750;
8'h0a : rvCrc[14] <= 32'h4c279971;
8'h0b : rvCrc[14] <= 32'h91287803;
8'h0c : rvCrc[14] <= 32'h8b85e533;
8'h0d : rvCrc[14] <= 32'h568a0441;
8'h0e : rvCrc[14] <= 32'h355b3a60;
8'h0f : rvCrc[14] <= 32'he854db12;
8'h10 : rvCrc[14] <= 32'he13391f3;
8'h11 : rvCrc[14] <= 32'h3c3c7081;
8'h12 : rvCrc[14] <= 32'h5fed4ea0;
8'h13 : rvCrc[14] <= 32'h82e2afd2;
8'h14 : rvCrc[14] <= 32'h984f32e2;
8'h15 : rvCrc[14] <= 32'h4540d390;
8'h16 : rvCrc[14] <= 32'h2691edb1;
8'h17 : rvCrc[14] <= 32'hfb9e0cc3;
8'h18 : rvCrc[14] <= 32'h13cad7d1;
8'h19 : rvCrc[14] <= 32'hcec536a3;
8'h1a : rvCrc[14] <= 32'had140882;
8'h1b : rvCrc[14] <= 32'h701be9f0;
8'h1c : rvCrc[14] <= 32'h6ab674c0;
8'h1d : rvCrc[14] <= 32'hb7b995b2;
8'h1e : rvCrc[14] <= 32'hd468ab93;
8'h1f : rvCrc[14] <= 32'h09674ae1;
8'h20 : rvCrc[14] <= 32'hc6a63e51;
8'h21 : rvCrc[14] <= 32'h1ba9df23;
8'h22 : rvCrc[14] <= 32'h7878e102;
8'h23 : rvCrc[14] <= 32'ha5770070;
8'h24 : rvCrc[14] <= 32'hbfda9d40;
8'h25 : rvCrc[14] <= 32'h62d57c32;
8'h26 : rvCrc[14] <= 32'h01044213;
8'h27 : rvCrc[14] <= 32'hdc0ba361;
8'h28 : rvCrc[14] <= 32'h345f7873;
8'h29 : rvCrc[14] <= 32'he9509901;
8'h2a : rvCrc[14] <= 32'h8a81a720;
8'h2b : rvCrc[14] <= 32'h578e4652;
8'h2c : rvCrc[14] <= 32'h4d23db62;
8'h2d : rvCrc[14] <= 32'h902c3a10;
8'h2e : rvCrc[14] <= 32'hf3fd0431;
8'h2f : rvCrc[14] <= 32'h2ef2e543;
8'h30 : rvCrc[14] <= 32'h2795afa2;
8'h31 : rvCrc[14] <= 32'hfa9a4ed0;
8'h32 : rvCrc[14] <= 32'h994b70f1;
8'h33 : rvCrc[14] <= 32'h44449183;
8'h34 : rvCrc[14] <= 32'h5ee90cb3;
8'h35 : rvCrc[14] <= 32'h83e6edc1;
8'h36 : rvCrc[14] <= 32'he037d3e0;
8'h37 : rvCrc[14] <= 32'h3d383292;
8'h38 : rvCrc[14] <= 32'hd56ce980;
8'h39 : rvCrc[14] <= 32'h086308f2;
8'h3a : rvCrc[14] <= 32'h6bb236d3;
8'h3b : rvCrc[14] <= 32'hb6bdd7a1;
8'h3c : rvCrc[14] <= 32'hac104a91;
8'h3d : rvCrc[14] <= 32'h711fabe3;
8'h3e : rvCrc[14] <= 32'h12ce95c2;
8'h3f : rvCrc[14] <= 32'hcfc174b0;
8'h40 : rvCrc[14] <= 32'h898d6115;
8'h41 : rvCrc[14] <= 32'h54828067;
8'h42 : rvCrc[14] <= 32'h3753be46;
8'h43 : rvCrc[14] <= 32'hea5c5f34;
8'h44 : rvCrc[14] <= 32'hf0f1c204;
8'h45 : rvCrc[14] <= 32'h2dfe2376;
8'h46 : rvCrc[14] <= 32'h4e2f1d57;
8'h47 : rvCrc[14] <= 32'h9320fc25;
8'h48 : rvCrc[14] <= 32'h7b742737;
8'h49 : rvCrc[14] <= 32'ha67bc645;
8'h4a : rvCrc[14] <= 32'hc5aaf864;
8'h4b : rvCrc[14] <= 32'h18a51916;
8'h4c : rvCrc[14] <= 32'h02088426;
8'h4d : rvCrc[14] <= 32'hdf076554;
8'h4e : rvCrc[14] <= 32'hbcd65b75;
8'h4f : rvCrc[14] <= 32'h61d9ba07;
8'h50 : rvCrc[14] <= 32'h68bef0e6;
8'h51 : rvCrc[14] <= 32'hb5b11194;
8'h52 : rvCrc[14] <= 32'hd6602fb5;
8'h53 : rvCrc[14] <= 32'h0b6fcec7;
8'h54 : rvCrc[14] <= 32'h11c253f7;
8'h55 : rvCrc[14] <= 32'hcccdb285;
8'h56 : rvCrc[14] <= 32'haf1c8ca4;
8'h57 : rvCrc[14] <= 32'h72136dd6;
8'h58 : rvCrc[14] <= 32'h9a47b6c4;
8'h59 : rvCrc[14] <= 32'h474857b6;
8'h5a : rvCrc[14] <= 32'h24996997;
8'h5b : rvCrc[14] <= 32'hf99688e5;
8'h5c : rvCrc[14] <= 32'he33b15d5;
8'h5d : rvCrc[14] <= 32'h3e34f4a7;
8'h5e : rvCrc[14] <= 32'h5de5ca86;
8'h5f : rvCrc[14] <= 32'h80ea2bf4;
8'h60 : rvCrc[14] <= 32'h4f2b5f44;
8'h61 : rvCrc[14] <= 32'h9224be36;
8'h62 : rvCrc[14] <= 32'hf1f58017;
8'h63 : rvCrc[14] <= 32'h2cfa6165;
8'h64 : rvCrc[14] <= 32'h3657fc55;
8'h65 : rvCrc[14] <= 32'heb581d27;
8'h66 : rvCrc[14] <= 32'h88892306;
8'h67 : rvCrc[14] <= 32'h5586c274;
8'h68 : rvCrc[14] <= 32'hbdd21966;
8'h69 : rvCrc[14] <= 32'h60ddf814;
8'h6a : rvCrc[14] <= 32'h030cc635;
8'h6b : rvCrc[14] <= 32'hde032747;
8'h6c : rvCrc[14] <= 32'hc4aeba77;
8'h6d : rvCrc[14] <= 32'h19a15b05;
8'h6e : rvCrc[14] <= 32'h7a706524;
8'h6f : rvCrc[14] <= 32'ha77f8456;
8'h70 : rvCrc[14] <= 32'hae18ceb7;
8'h71 : rvCrc[14] <= 32'h73172fc5;
8'h72 : rvCrc[14] <= 32'h10c611e4;
8'h73 : rvCrc[14] <= 32'hcdc9f096;
8'h74 : rvCrc[14] <= 32'hd7646da6;
8'h75 : rvCrc[14] <= 32'h0a6b8cd4;
8'h76 : rvCrc[14] <= 32'h69bab2f5;
8'h77 : rvCrc[14] <= 32'hb4b55387;
8'h78 : rvCrc[14] <= 32'h5ce18895;
8'h79 : rvCrc[14] <= 32'h81ee69e7;
8'h7a : rvCrc[14] <= 32'he23f57c6;
8'h7b : rvCrc[14] <= 32'h3f30b6b4;
8'h7c : rvCrc[14] <= 32'h259d2b84;
8'h7d : rvCrc[14] <= 32'hf892caf6;
8'h7e : rvCrc[14] <= 32'h9b43f4d7;
8'h7f : rvCrc[14] <= 32'h464c15a5;
8'h80 : rvCrc[14] <= 32'h17dbdf9d;
8'h81 : rvCrc[14] <= 32'hcad43eef;
8'h82 : rvCrc[14] <= 32'ha90500ce;
8'h83 : rvCrc[14] <= 32'h740ae1bc;
8'h84 : rvCrc[14] <= 32'h6ea77c8c;
8'h85 : rvCrc[14] <= 32'hb3a89dfe;
8'h86 : rvCrc[14] <= 32'hd079a3df;
8'h87 : rvCrc[14] <= 32'h0d7642ad;
8'h88 : rvCrc[14] <= 32'he52299bf;
8'h89 : rvCrc[14] <= 32'h382d78cd;
8'h8a : rvCrc[14] <= 32'h5bfc46ec;
8'h8b : rvCrc[14] <= 32'h86f3a79e;
8'h8c : rvCrc[14] <= 32'h9c5e3aae;
8'h8d : rvCrc[14] <= 32'h4151dbdc;
8'h8e : rvCrc[14] <= 32'h2280e5fd;
8'h8f : rvCrc[14] <= 32'hff8f048f;
8'h90 : rvCrc[14] <= 32'hf6e84e6e;
8'h91 : rvCrc[14] <= 32'h2be7af1c;
8'h92 : rvCrc[14] <= 32'h4836913d;
8'h93 : rvCrc[14] <= 32'h9539704f;
8'h94 : rvCrc[14] <= 32'h8f94ed7f;
8'h95 : rvCrc[14] <= 32'h529b0c0d;
8'h96 : rvCrc[14] <= 32'h314a322c;
8'h97 : rvCrc[14] <= 32'hec45d35e;
8'h98 : rvCrc[14] <= 32'h0411084c;
8'h99 : rvCrc[14] <= 32'hd91ee93e;
8'h9a : rvCrc[14] <= 32'hbacfd71f;
8'h9b : rvCrc[14] <= 32'h67c0366d;
8'h9c : rvCrc[14] <= 32'h7d6dab5d;
8'h9d : rvCrc[14] <= 32'ha0624a2f;
8'h9e : rvCrc[14] <= 32'hc3b3740e;
8'h9f : rvCrc[14] <= 32'h1ebc957c;
8'ha0 : rvCrc[14] <= 32'hd17de1cc;
8'ha1 : rvCrc[14] <= 32'h0c7200be;
8'ha2 : rvCrc[14] <= 32'h6fa33e9f;
8'ha3 : rvCrc[14] <= 32'hb2acdfed;
8'ha4 : rvCrc[14] <= 32'ha80142dd;
8'ha5 : rvCrc[14] <= 32'h750ea3af;
8'ha6 : rvCrc[14] <= 32'h16df9d8e;
8'ha7 : rvCrc[14] <= 32'hcbd07cfc;
8'ha8 : rvCrc[14] <= 32'h2384a7ee;
8'ha9 : rvCrc[14] <= 32'hfe8b469c;
8'haa : rvCrc[14] <= 32'h9d5a78bd;
8'hab : rvCrc[14] <= 32'h405599cf;
8'hac : rvCrc[14] <= 32'h5af804ff;
8'had : rvCrc[14] <= 32'h87f7e58d;
8'hae : rvCrc[14] <= 32'he426dbac;
8'haf : rvCrc[14] <= 32'h39293ade;
8'hb0 : rvCrc[14] <= 32'h304e703f;
8'hb1 : rvCrc[14] <= 32'hed41914d;
8'hb2 : rvCrc[14] <= 32'h8e90af6c;
8'hb3 : rvCrc[14] <= 32'h539f4e1e;
8'hb4 : rvCrc[14] <= 32'h4932d32e;
8'hb5 : rvCrc[14] <= 32'h943d325c;
8'hb6 : rvCrc[14] <= 32'hf7ec0c7d;
8'hb7 : rvCrc[14] <= 32'h2ae3ed0f;
8'hb8 : rvCrc[14] <= 32'hc2b7361d;
8'hb9 : rvCrc[14] <= 32'h1fb8d76f;
8'hba : rvCrc[14] <= 32'h7c69e94e;
8'hbb : rvCrc[14] <= 32'ha166083c;
8'hbc : rvCrc[14] <= 32'hbbcb950c;
8'hbd : rvCrc[14] <= 32'h66c4747e;
8'hbe : rvCrc[14] <= 32'h05154a5f;
8'hbf : rvCrc[14] <= 32'hd81aab2d;
8'hc0 : rvCrc[14] <= 32'h9e56be88;
8'hc1 : rvCrc[14] <= 32'h43595ffa;
8'hc2 : rvCrc[14] <= 32'h208861db;
8'hc3 : rvCrc[14] <= 32'hfd8780a9;
8'hc4 : rvCrc[14] <= 32'he72a1d99;
8'hc5 : rvCrc[14] <= 32'h3a25fceb;
8'hc6 : rvCrc[14] <= 32'h59f4c2ca;
8'hc7 : rvCrc[14] <= 32'h84fb23b8;
8'hc8 : rvCrc[14] <= 32'h6caff8aa;
8'hc9 : rvCrc[14] <= 32'hb1a019d8;
8'hca : rvCrc[14] <= 32'hd27127f9;
8'hcb : rvCrc[14] <= 32'h0f7ec68b;
8'hcc : rvCrc[14] <= 32'h15d35bbb;
8'hcd : rvCrc[14] <= 32'hc8dcbac9;
8'hce : rvCrc[14] <= 32'hab0d84e8;
8'hcf : rvCrc[14] <= 32'h7602659a;
8'hd0 : rvCrc[14] <= 32'h7f652f7b;
8'hd1 : rvCrc[14] <= 32'ha26ace09;
8'hd2 : rvCrc[14] <= 32'hc1bbf028;
8'hd3 : rvCrc[14] <= 32'h1cb4115a;
8'hd4 : rvCrc[14] <= 32'h06198c6a;
8'hd5 : rvCrc[14] <= 32'hdb166d18;
8'hd6 : rvCrc[14] <= 32'hb8c75339;
8'hd7 : rvCrc[14] <= 32'h65c8b24b;
8'hd8 : rvCrc[14] <= 32'h8d9c6959;
8'hd9 : rvCrc[14] <= 32'h5093882b;
8'hda : rvCrc[14] <= 32'h3342b60a;
8'hdb : rvCrc[14] <= 32'hee4d5778;
8'hdc : rvCrc[14] <= 32'hf4e0ca48;
8'hdd : rvCrc[14] <= 32'h29ef2b3a;
8'hde : rvCrc[14] <= 32'h4a3e151b;
8'hdf : rvCrc[14] <= 32'h9731f469;
8'he0 : rvCrc[14] <= 32'h58f080d9;
8'he1 : rvCrc[14] <= 32'h85ff61ab;
8'he2 : rvCrc[14] <= 32'he62e5f8a;
8'he3 : rvCrc[14] <= 32'h3b21bef8;
8'he4 : rvCrc[14] <= 32'h218c23c8;
8'he5 : rvCrc[14] <= 32'hfc83c2ba;
8'he6 : rvCrc[14] <= 32'h9f52fc9b;
8'he7 : rvCrc[14] <= 32'h425d1de9;
8'he8 : rvCrc[14] <= 32'haa09c6fb;
8'he9 : rvCrc[14] <= 32'h77062789;
8'hea : rvCrc[14] <= 32'h14d719a8;
8'heb : rvCrc[14] <= 32'hc9d8f8da;
8'hec : rvCrc[14] <= 32'hd37565ea;
8'hed : rvCrc[14] <= 32'h0e7a8498;
8'hee : rvCrc[14] <= 32'h6dabbab9;
8'hef : rvCrc[14] <= 32'hb0a45bcb;
8'hf0 : rvCrc[14] <= 32'hb9c3112a;
8'hf1 : rvCrc[14] <= 32'h64ccf058;
8'hf2 : rvCrc[14] <= 32'h071dce79;
8'hf3 : rvCrc[14] <= 32'hda122f0b;
8'hf4 : rvCrc[14] <= 32'hc0bfb23b;
8'hf5 : rvCrc[14] <= 32'h1db05349;
8'hf6 : rvCrc[14] <= 32'h7e616d68;
8'hf7 : rvCrc[14] <= 32'ha36e8c1a;
8'hf8 : rvCrc[14] <= 32'h4b3a5708;
8'hf9 : rvCrc[14] <= 32'h9635b67a;
8'hfa : rvCrc[14] <= 32'hf5e4885b;
8'hfb : rvCrc[14] <= 32'h28eb6929;
8'hfc : rvCrc[14] <= 32'h3246f419;
8'hfd : rvCrc[14] <= 32'hef49156b;
8'hfe : rvCrc[14] <= 32'h8c982b4a;
8'hff : rvCrc[14] <= 32'h5197ca38;
endcase
case(iv_Input[127:120])
8'h00 : rvCrc[15] <= 32'h00000000;
8'h01 : rvCrc[15] <= 32'h2fb7bf3a;
8'h02 : rvCrc[15] <= 32'h5f6f7e74;
8'h03 : rvCrc[15] <= 32'h70d8c14e;
8'h04 : rvCrc[15] <= 32'hbedefce8;
8'h05 : rvCrc[15] <= 32'h916943d2;
8'h06 : rvCrc[15] <= 32'he1b1829c;
8'h07 : rvCrc[15] <= 32'hce063da6;
8'h08 : rvCrc[15] <= 32'h797ce467;
8'h09 : rvCrc[15] <= 32'h56cb5b5d;
8'h0a : rvCrc[15] <= 32'h26139a13;
8'h0b : rvCrc[15] <= 32'h09a42529;
8'h0c : rvCrc[15] <= 32'hc7a2188f;
8'h0d : rvCrc[15] <= 32'he815a7b5;
8'h0e : rvCrc[15] <= 32'h98cd66fb;
8'h0f : rvCrc[15] <= 32'hb77ad9c1;
8'h10 : rvCrc[15] <= 32'hf2f9c8ce;
8'h11 : rvCrc[15] <= 32'hdd4e77f4;
8'h12 : rvCrc[15] <= 32'had96b6ba;
8'h13 : rvCrc[15] <= 32'h82210980;
8'h14 : rvCrc[15] <= 32'h4c273426;
8'h15 : rvCrc[15] <= 32'h63908b1c;
8'h16 : rvCrc[15] <= 32'h13484a52;
8'h17 : rvCrc[15] <= 32'h3cfff568;
8'h18 : rvCrc[15] <= 32'h8b852ca9;
8'h19 : rvCrc[15] <= 32'ha4329393;
8'h1a : rvCrc[15] <= 32'hd4ea52dd;
8'h1b : rvCrc[15] <= 32'hfb5dede7;
8'h1c : rvCrc[15] <= 32'h355bd041;
8'h1d : rvCrc[15] <= 32'h1aec6f7b;
8'h1e : rvCrc[15] <= 32'h6a34ae35;
8'h1f : rvCrc[15] <= 32'h4583110f;
8'h20 : rvCrc[15] <= 32'he1328c2b;
8'h21 : rvCrc[15] <= 32'hce853311;
8'h22 : rvCrc[15] <= 32'hbe5df25f;
8'h23 : rvCrc[15] <= 32'h91ea4d65;
8'h24 : rvCrc[15] <= 32'h5fec70c3;
8'h25 : rvCrc[15] <= 32'h705bcff9;
8'h26 : rvCrc[15] <= 32'h00830eb7;
8'h27 : rvCrc[15] <= 32'h2f34b18d;
8'h28 : rvCrc[15] <= 32'h984e684c;
8'h29 : rvCrc[15] <= 32'hb7f9d776;
8'h2a : rvCrc[15] <= 32'hc7211638;
8'h2b : rvCrc[15] <= 32'he896a902;
8'h2c : rvCrc[15] <= 32'h269094a4;
8'h2d : rvCrc[15] <= 32'h09272b9e;
8'h2e : rvCrc[15] <= 32'h79ffead0;
8'h2f : rvCrc[15] <= 32'h564855ea;
8'h30 : rvCrc[15] <= 32'h13cb44e5;
8'h31 : rvCrc[15] <= 32'h3c7cfbdf;
8'h32 : rvCrc[15] <= 32'h4ca43a91;
8'h33 : rvCrc[15] <= 32'h631385ab;
8'h34 : rvCrc[15] <= 32'had15b80d;
8'h35 : rvCrc[15] <= 32'h82a20737;
8'h36 : rvCrc[15] <= 32'hf27ac679;
8'h37 : rvCrc[15] <= 32'hddcd7943;
8'h38 : rvCrc[15] <= 32'h6ab7a082;
8'h39 : rvCrc[15] <= 32'h45001fb8;
8'h3a : rvCrc[15] <= 32'h35d8def6;
8'h3b : rvCrc[15] <= 32'h1a6f61cc;
8'h3c : rvCrc[15] <= 32'hd4695c6a;
8'h3d : rvCrc[15] <= 32'hfbdee350;
8'h3e : rvCrc[15] <= 32'h8b06221e;
8'h3f : rvCrc[15] <= 32'ha4b19d24;
8'h40 : rvCrc[15] <= 32'hc6a405e1;
8'h41 : rvCrc[15] <= 32'he913badb;
8'h42 : rvCrc[15] <= 32'h99cb7b95;
8'h43 : rvCrc[15] <= 32'hb67cc4af;
8'h44 : rvCrc[15] <= 32'h787af909;
8'h45 : rvCrc[15] <= 32'h57cd4633;
8'h46 : rvCrc[15] <= 32'h2715877d;
8'h47 : rvCrc[15] <= 32'h08a23847;
8'h48 : rvCrc[15] <= 32'hbfd8e186;
8'h49 : rvCrc[15] <= 32'h906f5ebc;
8'h4a : rvCrc[15] <= 32'he0b79ff2;
8'h4b : rvCrc[15] <= 32'hcf0020c8;
8'h4c : rvCrc[15] <= 32'h01061d6e;
8'h4d : rvCrc[15] <= 32'h2eb1a254;
8'h4e : rvCrc[15] <= 32'h5e69631a;
8'h4f : rvCrc[15] <= 32'h71dedc20;
8'h50 : rvCrc[15] <= 32'h345dcd2f;
8'h51 : rvCrc[15] <= 32'h1bea7215;
8'h52 : rvCrc[15] <= 32'h6b32b35b;
8'h53 : rvCrc[15] <= 32'h44850c61;
8'h54 : rvCrc[15] <= 32'h8a8331c7;
8'h55 : rvCrc[15] <= 32'ha5348efd;
8'h56 : rvCrc[15] <= 32'hd5ec4fb3;
8'h57 : rvCrc[15] <= 32'hfa5bf089;
8'h58 : rvCrc[15] <= 32'h4d212948;
8'h59 : rvCrc[15] <= 32'h62969672;
8'h5a : rvCrc[15] <= 32'h124e573c;
8'h5b : rvCrc[15] <= 32'h3df9e806;
8'h5c : rvCrc[15] <= 32'hf3ffd5a0;
8'h5d : rvCrc[15] <= 32'hdc486a9a;
8'h5e : rvCrc[15] <= 32'hac90abd4;
8'h5f : rvCrc[15] <= 32'h832714ee;
8'h60 : rvCrc[15] <= 32'h279689ca;
8'h61 : rvCrc[15] <= 32'h082136f0;
8'h62 : rvCrc[15] <= 32'h78f9f7be;
8'h63 : rvCrc[15] <= 32'h574e4884;
8'h64 : rvCrc[15] <= 32'h99487522;
8'h65 : rvCrc[15] <= 32'hb6ffca18;
8'h66 : rvCrc[15] <= 32'hc6270b56;
8'h67 : rvCrc[15] <= 32'he990b46c;
8'h68 : rvCrc[15] <= 32'h5eea6dad;
8'h69 : rvCrc[15] <= 32'h715dd297;
8'h6a : rvCrc[15] <= 32'h018513d9;
8'h6b : rvCrc[15] <= 32'h2e32ace3;
8'h6c : rvCrc[15] <= 32'he0349145;
8'h6d : rvCrc[15] <= 32'hcf832e7f;
8'h6e : rvCrc[15] <= 32'hbf5bef31;
8'h6f : rvCrc[15] <= 32'h90ec500b;
8'h70 : rvCrc[15] <= 32'hd56f4104;
8'h71 : rvCrc[15] <= 32'hfad8fe3e;
8'h72 : rvCrc[15] <= 32'h8a003f70;
8'h73 : rvCrc[15] <= 32'ha5b7804a;
8'h74 : rvCrc[15] <= 32'h6bb1bdec;
8'h75 : rvCrc[15] <= 32'h440602d6;
8'h76 : rvCrc[15] <= 32'h34dec398;
8'h77 : rvCrc[15] <= 32'h1b697ca2;
8'h78 : rvCrc[15] <= 32'hac13a563;
8'h79 : rvCrc[15] <= 32'h83a41a59;
8'h7a : rvCrc[15] <= 32'hf37cdb17;
8'h7b : rvCrc[15] <= 32'hdccb642d;
8'h7c : rvCrc[15] <= 32'h12cd598b;
8'h7d : rvCrc[15] <= 32'h3d7ae6b1;
8'h7e : rvCrc[15] <= 32'h4da227ff;
8'h7f : rvCrc[15] <= 32'h621598c5;
8'h80 : rvCrc[15] <= 32'h89891675;
8'h81 : rvCrc[15] <= 32'ha63ea94f;
8'h82 : rvCrc[15] <= 32'hd6e66801;
8'h83 : rvCrc[15] <= 32'hf951d73b;
8'h84 : rvCrc[15] <= 32'h3757ea9d;
8'h85 : rvCrc[15] <= 32'h18e055a7;
8'h86 : rvCrc[15] <= 32'h683894e9;
8'h87 : rvCrc[15] <= 32'h478f2bd3;
8'h88 : rvCrc[15] <= 32'hf0f5f212;
8'h89 : rvCrc[15] <= 32'hdf424d28;
8'h8a : rvCrc[15] <= 32'haf9a8c66;
8'h8b : rvCrc[15] <= 32'h802d335c;
8'h8c : rvCrc[15] <= 32'h4e2b0efa;
8'h8d : rvCrc[15] <= 32'h619cb1c0;
8'h8e : rvCrc[15] <= 32'h1144708e;
8'h8f : rvCrc[15] <= 32'h3ef3cfb4;
8'h90 : rvCrc[15] <= 32'h7b70debb;
8'h91 : rvCrc[15] <= 32'h54c76181;
8'h92 : rvCrc[15] <= 32'h241fa0cf;
8'h93 : rvCrc[15] <= 32'h0ba81ff5;
8'h94 : rvCrc[15] <= 32'hc5ae2253;
8'h95 : rvCrc[15] <= 32'hea199d69;
8'h96 : rvCrc[15] <= 32'h9ac15c27;
8'h97 : rvCrc[15] <= 32'hb576e31d;
8'h98 : rvCrc[15] <= 32'h020c3adc;
8'h99 : rvCrc[15] <= 32'h2dbb85e6;
8'h9a : rvCrc[15] <= 32'h5d6344a8;
8'h9b : rvCrc[15] <= 32'h72d4fb92;
8'h9c : rvCrc[15] <= 32'hbcd2c634;
8'h9d : rvCrc[15] <= 32'h9365790e;
8'h9e : rvCrc[15] <= 32'he3bdb840;
8'h9f : rvCrc[15] <= 32'hcc0a077a;
8'ha0 : rvCrc[15] <= 32'h68bb9a5e;
8'ha1 : rvCrc[15] <= 32'h470c2564;
8'ha2 : rvCrc[15] <= 32'h37d4e42a;
8'ha3 : rvCrc[15] <= 32'h18635b10;
8'ha4 : rvCrc[15] <= 32'hd66566b6;
8'ha5 : rvCrc[15] <= 32'hf9d2d98c;
8'ha6 : rvCrc[15] <= 32'h890a18c2;
8'ha7 : rvCrc[15] <= 32'ha6bda7f8;
8'ha8 : rvCrc[15] <= 32'h11c77e39;
8'ha9 : rvCrc[15] <= 32'h3e70c103;
8'haa : rvCrc[15] <= 32'h4ea8004d;
8'hab : rvCrc[15] <= 32'h611fbf77;
8'hac : rvCrc[15] <= 32'haf1982d1;
8'had : rvCrc[15] <= 32'h80ae3deb;
8'hae : rvCrc[15] <= 32'hf076fca5;
8'haf : rvCrc[15] <= 32'hdfc1439f;
8'hb0 : rvCrc[15] <= 32'h9a425290;
8'hb1 : rvCrc[15] <= 32'hb5f5edaa;
8'hb2 : rvCrc[15] <= 32'hc52d2ce4;
8'hb3 : rvCrc[15] <= 32'hea9a93de;
8'hb4 : rvCrc[15] <= 32'h249cae78;
8'hb5 : rvCrc[15] <= 32'h0b2b1142;
8'hb6 : rvCrc[15] <= 32'h7bf3d00c;
8'hb7 : rvCrc[15] <= 32'h54446f36;
8'hb8 : rvCrc[15] <= 32'he33eb6f7;
8'hb9 : rvCrc[15] <= 32'hcc8909cd;
8'hba : rvCrc[15] <= 32'hbc51c883;
8'hbb : rvCrc[15] <= 32'h93e677b9;
8'hbc : rvCrc[15] <= 32'h5de04a1f;
8'hbd : rvCrc[15] <= 32'h7257f525;
8'hbe : rvCrc[15] <= 32'h028f346b;
8'hbf : rvCrc[15] <= 32'h2d388b51;
8'hc0 : rvCrc[15] <= 32'h4f2d1394;
8'hc1 : rvCrc[15] <= 32'h609aacae;
8'hc2 : rvCrc[15] <= 32'h10426de0;
8'hc3 : rvCrc[15] <= 32'h3ff5d2da;
8'hc4 : rvCrc[15] <= 32'hf1f3ef7c;
8'hc5 : rvCrc[15] <= 32'hde445046;
8'hc6 : rvCrc[15] <= 32'hae9c9108;
8'hc7 : rvCrc[15] <= 32'h812b2e32;
8'hc8 : rvCrc[15] <= 32'h3651f7f3;
8'hc9 : rvCrc[15] <= 32'h19e648c9;
8'hca : rvCrc[15] <= 32'h693e8987;
8'hcb : rvCrc[15] <= 32'h468936bd;
8'hcc : rvCrc[15] <= 32'h888f0b1b;
8'hcd : rvCrc[15] <= 32'ha738b421;
8'hce : rvCrc[15] <= 32'hd7e0756f;
8'hcf : rvCrc[15] <= 32'hf857ca55;
8'hd0 : rvCrc[15] <= 32'hbdd4db5a;
8'hd1 : rvCrc[15] <= 32'h92636460;
8'hd2 : rvCrc[15] <= 32'he2bba52e;
8'hd3 : rvCrc[15] <= 32'hcd0c1a14;
8'hd4 : rvCrc[15] <= 32'h030a27b2;
8'hd5 : rvCrc[15] <= 32'h2cbd9888;
8'hd6 : rvCrc[15] <= 32'h5c6559c6;
8'hd7 : rvCrc[15] <= 32'h73d2e6fc;
8'hd8 : rvCrc[15] <= 32'hc4a83f3d;
8'hd9 : rvCrc[15] <= 32'heb1f8007;
8'hda : rvCrc[15] <= 32'h9bc74149;
8'hdb : rvCrc[15] <= 32'hb470fe73;
8'hdc : rvCrc[15] <= 32'h7a76c3d5;
8'hdd : rvCrc[15] <= 32'h55c17cef;
8'hde : rvCrc[15] <= 32'h2519bda1;
8'hdf : rvCrc[15] <= 32'h0aae029b;
8'he0 : rvCrc[15] <= 32'hae1f9fbf;
8'he1 : rvCrc[15] <= 32'h81a82085;
8'he2 : rvCrc[15] <= 32'hf170e1cb;
8'he3 : rvCrc[15] <= 32'hdec75ef1;
8'he4 : rvCrc[15] <= 32'h10c16357;
8'he5 : rvCrc[15] <= 32'h3f76dc6d;
8'he6 : rvCrc[15] <= 32'h4fae1d23;
8'he7 : rvCrc[15] <= 32'h6019a219;
8'he8 : rvCrc[15] <= 32'hd7637bd8;
8'he9 : rvCrc[15] <= 32'hf8d4c4e2;
8'hea : rvCrc[15] <= 32'h880c05ac;
8'heb : rvCrc[15] <= 32'ha7bbba96;
8'hec : rvCrc[15] <= 32'h69bd8730;
8'hed : rvCrc[15] <= 32'h460a380a;
8'hee : rvCrc[15] <= 32'h36d2f944;
8'hef : rvCrc[15] <= 32'h1965467e;
8'hf0 : rvCrc[15] <= 32'h5ce65771;
8'hf1 : rvCrc[15] <= 32'h7351e84b;
8'hf2 : rvCrc[15] <= 32'h03892905;
8'hf3 : rvCrc[15] <= 32'h2c3e963f;
8'hf4 : rvCrc[15] <= 32'he238ab99;
8'hf5 : rvCrc[15] <= 32'hcd8f14a3;
8'hf6 : rvCrc[15] <= 32'hbd57d5ed;
8'hf7 : rvCrc[15] <= 32'h92e06ad7;
8'hf8 : rvCrc[15] <= 32'h259ab316;
8'hf9 : rvCrc[15] <= 32'h0a2d0c2c;
8'hfa : rvCrc[15] <= 32'h7af5cd62;
8'hfb : rvCrc[15] <= 32'h55427258;
8'hfc : rvCrc[15] <= 32'h9b444ffe;
8'hfd : rvCrc[15] <= 32'hb4f3f0c4;
8'hfe : rvCrc[15] <= 32'hc42b318a;
8'hff : rvCrc[15] <= 32'heb9c8eb0;
endcase
case(iv_Input[135:128])
8'h00 : rvCrc[16] <= 32'h00000000;
8'h01 : rvCrc[16] <= 32'h17d3315d;
8'h02 : rvCrc[16] <= 32'h2fa662ba;
8'h03 : rvCrc[16] <= 32'h387553e7;
8'h04 : rvCrc[16] <= 32'h5f4cc574;
8'h05 : rvCrc[16] <= 32'h489ff429;
8'h06 : rvCrc[16] <= 32'h70eaa7ce;
8'h07 : rvCrc[16] <= 32'h67399693;
8'h08 : rvCrc[16] <= 32'hbe998ae8;
8'h09 : rvCrc[16] <= 32'ha94abbb5;
8'h0a : rvCrc[16] <= 32'h913fe852;
8'h0b : rvCrc[16] <= 32'h86ecd90f;
8'h0c : rvCrc[16] <= 32'he1d54f9c;
8'h0d : rvCrc[16] <= 32'hf6067ec1;
8'h0e : rvCrc[16] <= 32'hce732d26;
8'h0f : rvCrc[16] <= 32'hd9a01c7b;
8'h10 : rvCrc[16] <= 32'h79f20867;
8'h11 : rvCrc[16] <= 32'h6e21393a;
8'h12 : rvCrc[16] <= 32'h56546add;
8'h13 : rvCrc[16] <= 32'h41875b80;
8'h14 : rvCrc[16] <= 32'h26becd13;
8'h15 : rvCrc[16] <= 32'h316dfc4e;
8'h16 : rvCrc[16] <= 32'h0918afa9;
8'h17 : rvCrc[16] <= 32'h1ecb9ef4;
8'h18 : rvCrc[16] <= 32'hc76b828f;
8'h19 : rvCrc[16] <= 32'hd0b8b3d2;
8'h1a : rvCrc[16] <= 32'he8cde035;
8'h1b : rvCrc[16] <= 32'hff1ed168;
8'h1c : rvCrc[16] <= 32'h982747fb;
8'h1d : rvCrc[16] <= 32'h8ff476a6;
8'h1e : rvCrc[16] <= 32'hb7812541;
8'h1f : rvCrc[16] <= 32'ha052141c;
8'h20 : rvCrc[16] <= 32'hf3e410ce;
8'h21 : rvCrc[16] <= 32'he4372193;
8'h22 : rvCrc[16] <= 32'hdc427274;
8'h23 : rvCrc[16] <= 32'hcb914329;
8'h24 : rvCrc[16] <= 32'haca8d5ba;
8'h25 : rvCrc[16] <= 32'hbb7be4e7;
8'h26 : rvCrc[16] <= 32'h830eb700;
8'h27 : rvCrc[16] <= 32'h94dd865d;
8'h28 : rvCrc[16] <= 32'h4d7d9a26;
8'h29 : rvCrc[16] <= 32'h5aaeab7b;
8'h2a : rvCrc[16] <= 32'h62dbf89c;
8'h2b : rvCrc[16] <= 32'h7508c9c1;
8'h2c : rvCrc[16] <= 32'h12315f52;
8'h2d : rvCrc[16] <= 32'h05e26e0f;
8'h2e : rvCrc[16] <= 32'h3d973de8;
8'h2f : rvCrc[16] <= 32'h2a440cb5;
8'h30 : rvCrc[16] <= 32'h8a1618a9;
8'h31 : rvCrc[16] <= 32'h9dc529f4;
8'h32 : rvCrc[16] <= 32'ha5b07a13;
8'h33 : rvCrc[16] <= 32'hb2634b4e;
8'h34 : rvCrc[16] <= 32'hd55adddd;
8'h35 : rvCrc[16] <= 32'hc289ec80;
8'h36 : rvCrc[16] <= 32'hfafcbf67;
8'h37 : rvCrc[16] <= 32'hed2f8e3a;
8'h38 : rvCrc[16] <= 32'h348f9241;
8'h39 : rvCrc[16] <= 32'h235ca31c;
8'h3a : rvCrc[16] <= 32'h1b29f0fb;
8'h3b : rvCrc[16] <= 32'h0cfac1a6;
8'h3c : rvCrc[16] <= 32'h6bc35735;
8'h3d : rvCrc[16] <= 32'h7c106668;
8'h3e : rvCrc[16] <= 32'h4465358f;
8'h3f : rvCrc[16] <= 32'h53b604d2;
8'h40 : rvCrc[16] <= 32'he3093c2b;
8'h41 : rvCrc[16] <= 32'hf4da0d76;
8'h42 : rvCrc[16] <= 32'hccaf5e91;
8'h43 : rvCrc[16] <= 32'hdb7c6fcc;
8'h44 : rvCrc[16] <= 32'hbc45f95f;
8'h45 : rvCrc[16] <= 32'hab96c802;
8'h46 : rvCrc[16] <= 32'h93e39be5;
8'h47 : rvCrc[16] <= 32'h8430aab8;
8'h48 : rvCrc[16] <= 32'h5d90b6c3;
8'h49 : rvCrc[16] <= 32'h4a43879e;
8'h4a : rvCrc[16] <= 32'h7236d479;
8'h4b : rvCrc[16] <= 32'h65e5e524;
8'h4c : rvCrc[16] <= 32'h02dc73b7;
8'h4d : rvCrc[16] <= 32'h150f42ea;
8'h4e : rvCrc[16] <= 32'h2d7a110d;
8'h4f : rvCrc[16] <= 32'h3aa92050;
8'h50 : rvCrc[16] <= 32'h9afb344c;
8'h51 : rvCrc[16] <= 32'h8d280511;
8'h52 : rvCrc[16] <= 32'hb55d56f6;
8'h53 : rvCrc[16] <= 32'ha28e67ab;
8'h54 : rvCrc[16] <= 32'hc5b7f138;
8'h55 : rvCrc[16] <= 32'hd264c065;
8'h56 : rvCrc[16] <= 32'hea119382;
8'h57 : rvCrc[16] <= 32'hfdc2a2df;
8'h58 : rvCrc[16] <= 32'h2462bea4;
8'h59 : rvCrc[16] <= 32'h33b18ff9;
8'h5a : rvCrc[16] <= 32'h0bc4dc1e;
8'h5b : rvCrc[16] <= 32'h1c17ed43;
8'h5c : rvCrc[16] <= 32'h7b2e7bd0;
8'h5d : rvCrc[16] <= 32'h6cfd4a8d;
8'h5e : rvCrc[16] <= 32'h5488196a;
8'h5f : rvCrc[16] <= 32'h435b2837;
8'h60 : rvCrc[16] <= 32'h10ed2ce5;
8'h61 : rvCrc[16] <= 32'h073e1db8;
8'h62 : rvCrc[16] <= 32'h3f4b4e5f;
8'h63 : rvCrc[16] <= 32'h28987f02;
8'h64 : rvCrc[16] <= 32'h4fa1e991;
8'h65 : rvCrc[16] <= 32'h5872d8cc;
8'h66 : rvCrc[16] <= 32'h60078b2b;
8'h67 : rvCrc[16] <= 32'h77d4ba76;
8'h68 : rvCrc[16] <= 32'hae74a60d;
8'h69 : rvCrc[16] <= 32'hb9a79750;
8'h6a : rvCrc[16] <= 32'h81d2c4b7;
8'h6b : rvCrc[16] <= 32'h9601f5ea;
8'h6c : rvCrc[16] <= 32'hf1386379;
8'h6d : rvCrc[16] <= 32'he6eb5224;
8'h6e : rvCrc[16] <= 32'hde9e01c3;
8'h6f : rvCrc[16] <= 32'hc94d309e;
8'h70 : rvCrc[16] <= 32'h691f2482;
8'h71 : rvCrc[16] <= 32'h7ecc15df;
8'h72 : rvCrc[16] <= 32'h46b94638;
8'h73 : rvCrc[16] <= 32'h516a7765;
8'h74 : rvCrc[16] <= 32'h3653e1f6;
8'h75 : rvCrc[16] <= 32'h2180d0ab;
8'h76 : rvCrc[16] <= 32'h19f5834c;
8'h77 : rvCrc[16] <= 32'h0e26b211;
8'h78 : rvCrc[16] <= 32'hd786ae6a;
8'h79 : rvCrc[16] <= 32'hc0559f37;
8'h7a : rvCrc[16] <= 32'hf820ccd0;
8'h7b : rvCrc[16] <= 32'heff3fd8d;
8'h7c : rvCrc[16] <= 32'h88ca6b1e;
8'h7d : rvCrc[16] <= 32'h9f195a43;
8'h7e : rvCrc[16] <= 32'ha76c09a4;
8'h7f : rvCrc[16] <= 32'hb0bf38f9;
8'h80 : rvCrc[16] <= 32'hc2d365e1;
8'h81 : rvCrc[16] <= 32'hd50054bc;
8'h82 : rvCrc[16] <= 32'hed75075b;
8'h83 : rvCrc[16] <= 32'hfaa63606;
8'h84 : rvCrc[16] <= 32'h9d9fa095;
8'h85 : rvCrc[16] <= 32'h8a4c91c8;
8'h86 : rvCrc[16] <= 32'hb239c22f;
8'h87 : rvCrc[16] <= 32'ha5eaf372;
8'h88 : rvCrc[16] <= 32'h7c4aef09;
8'h89 : rvCrc[16] <= 32'h6b99de54;
8'h8a : rvCrc[16] <= 32'h53ec8db3;
8'h8b : rvCrc[16] <= 32'h443fbcee;
8'h8c : rvCrc[16] <= 32'h23062a7d;
8'h8d : rvCrc[16] <= 32'h34d51b20;
8'h8e : rvCrc[16] <= 32'h0ca048c7;
8'h8f : rvCrc[16] <= 32'h1b73799a;
8'h90 : rvCrc[16] <= 32'hbb216d86;
8'h91 : rvCrc[16] <= 32'hacf25cdb;
8'h92 : rvCrc[16] <= 32'h94870f3c;
8'h93 : rvCrc[16] <= 32'h83543e61;
8'h94 : rvCrc[16] <= 32'he46da8f2;
8'h95 : rvCrc[16] <= 32'hf3be99af;
8'h96 : rvCrc[16] <= 32'hcbcbca48;
8'h97 : rvCrc[16] <= 32'hdc18fb15;
8'h98 : rvCrc[16] <= 32'h05b8e76e;
8'h99 : rvCrc[16] <= 32'h126bd633;
8'h9a : rvCrc[16] <= 32'h2a1e85d4;
8'h9b : rvCrc[16] <= 32'h3dcdb489;
8'h9c : rvCrc[16] <= 32'h5af4221a;
8'h9d : rvCrc[16] <= 32'h4d271347;
8'h9e : rvCrc[16] <= 32'h755240a0;
8'h9f : rvCrc[16] <= 32'h628171fd;
8'ha0 : rvCrc[16] <= 32'h3137752f;
8'ha1 : rvCrc[16] <= 32'h26e44472;
8'ha2 : rvCrc[16] <= 32'h1e911795;
8'ha3 : rvCrc[16] <= 32'h094226c8;
8'ha4 : rvCrc[16] <= 32'h6e7bb05b;
8'ha5 : rvCrc[16] <= 32'h79a88106;
8'ha6 : rvCrc[16] <= 32'h41ddd2e1;
8'ha7 : rvCrc[16] <= 32'h560ee3bc;
8'ha8 : rvCrc[16] <= 32'h8faeffc7;
8'ha9 : rvCrc[16] <= 32'h987dce9a;
8'haa : rvCrc[16] <= 32'ha0089d7d;
8'hab : rvCrc[16] <= 32'hb7dbac20;
8'hac : rvCrc[16] <= 32'hd0e23ab3;
8'had : rvCrc[16] <= 32'hc7310bee;
8'hae : rvCrc[16] <= 32'hff445809;
8'haf : rvCrc[16] <= 32'he8976954;
8'hb0 : rvCrc[16] <= 32'h48c57d48;
8'hb1 : rvCrc[16] <= 32'h5f164c15;
8'hb2 : rvCrc[16] <= 32'h67631ff2;
8'hb3 : rvCrc[16] <= 32'h70b02eaf;
8'hb4 : rvCrc[16] <= 32'h1789b83c;
8'hb5 : rvCrc[16] <= 32'h005a8961;
8'hb6 : rvCrc[16] <= 32'h382fda86;
8'hb7 : rvCrc[16] <= 32'h2ffcebdb;
8'hb8 : rvCrc[16] <= 32'hf65cf7a0;
8'hb9 : rvCrc[16] <= 32'he18fc6fd;
8'hba : rvCrc[16] <= 32'hd9fa951a;
8'hbb : rvCrc[16] <= 32'hce29a447;
8'hbc : rvCrc[16] <= 32'ha91032d4;
8'hbd : rvCrc[16] <= 32'hbec30389;
8'hbe : rvCrc[16] <= 32'h86b6506e;
8'hbf : rvCrc[16] <= 32'h91656133;
8'hc0 : rvCrc[16] <= 32'h21da59ca;
8'hc1 : rvCrc[16] <= 32'h36096897;
8'hc2 : rvCrc[16] <= 32'h0e7c3b70;
8'hc3 : rvCrc[16] <= 32'h19af0a2d;
8'hc4 : rvCrc[16] <= 32'h7e969cbe;
8'hc5 : rvCrc[16] <= 32'h6945ade3;
8'hc6 : rvCrc[16] <= 32'h5130fe04;
8'hc7 : rvCrc[16] <= 32'h46e3cf59;
8'hc8 : rvCrc[16] <= 32'h9f43d322;
8'hc9 : rvCrc[16] <= 32'h8890e27f;
8'hca : rvCrc[16] <= 32'hb0e5b198;
8'hcb : rvCrc[16] <= 32'ha73680c5;
8'hcc : rvCrc[16] <= 32'hc00f1656;
8'hcd : rvCrc[16] <= 32'hd7dc270b;
8'hce : rvCrc[16] <= 32'hefa974ec;
8'hcf : rvCrc[16] <= 32'hf87a45b1;
8'hd0 : rvCrc[16] <= 32'h582851ad;
8'hd1 : rvCrc[16] <= 32'h4ffb60f0;
8'hd2 : rvCrc[16] <= 32'h778e3317;
8'hd3 : rvCrc[16] <= 32'h605d024a;
8'hd4 : rvCrc[16] <= 32'h076494d9;
8'hd5 : rvCrc[16] <= 32'h10b7a584;
8'hd6 : rvCrc[16] <= 32'h28c2f663;
8'hd7 : rvCrc[16] <= 32'h3f11c73e;
8'hd8 : rvCrc[16] <= 32'he6b1db45;
8'hd9 : rvCrc[16] <= 32'hf162ea18;
8'hda : rvCrc[16] <= 32'hc917b9ff;
8'hdb : rvCrc[16] <= 32'hdec488a2;
8'hdc : rvCrc[16] <= 32'hb9fd1e31;
8'hdd : rvCrc[16] <= 32'hae2e2f6c;
8'hde : rvCrc[16] <= 32'h965b7c8b;
8'hdf : rvCrc[16] <= 32'h81884dd6;
8'he0 : rvCrc[16] <= 32'hd23e4904;
8'he1 : rvCrc[16] <= 32'hc5ed7859;
8'he2 : rvCrc[16] <= 32'hfd982bbe;
8'he3 : rvCrc[16] <= 32'hea4b1ae3;
8'he4 : rvCrc[16] <= 32'h8d728c70;
8'he5 : rvCrc[16] <= 32'h9aa1bd2d;
8'he6 : rvCrc[16] <= 32'ha2d4eeca;
8'he7 : rvCrc[16] <= 32'hb507df97;
8'he8 : rvCrc[16] <= 32'h6ca7c3ec;
8'he9 : rvCrc[16] <= 32'h7b74f2b1;
8'hea : rvCrc[16] <= 32'h4301a156;
8'heb : rvCrc[16] <= 32'h54d2900b;
8'hec : rvCrc[16] <= 32'h33eb0698;
8'hed : rvCrc[16] <= 32'h243837c5;
8'hee : rvCrc[16] <= 32'h1c4d6422;
8'hef : rvCrc[16] <= 32'h0b9e557f;
8'hf0 : rvCrc[16] <= 32'habcc4163;
8'hf1 : rvCrc[16] <= 32'hbc1f703e;
8'hf2 : rvCrc[16] <= 32'h846a23d9;
8'hf3 : rvCrc[16] <= 32'h93b91284;
8'hf4 : rvCrc[16] <= 32'hf4808417;
8'hf5 : rvCrc[16] <= 32'he353b54a;
8'hf6 : rvCrc[16] <= 32'hdb26e6ad;
8'hf7 : rvCrc[16] <= 32'hccf5d7f0;
8'hf8 : rvCrc[16] <= 32'h1555cb8b;
8'hf9 : rvCrc[16] <= 32'h0286fad6;
8'hfa : rvCrc[16] <= 32'h3af3a931;
8'hfb : rvCrc[16] <= 32'h2d20986c;
8'hfc : rvCrc[16] <= 32'h4a190eff;
8'hfd : rvCrc[16] <= 32'h5dca3fa2;
8'hfe : rvCrc[16] <= 32'h65bf6c45;
8'hff : rvCrc[16] <= 32'h726c5d18;
endcase
case(iv_Input[143:136])
8'h00 : rvCrc[17] <= 32'h00000000;
8'h01 : rvCrc[17] <= 32'h8167d675;
8'h02 : rvCrc[17] <= 32'h060eb15d;
8'h03 : rvCrc[17] <= 32'h87696728;
8'h04 : rvCrc[17] <= 32'h0c1d62ba;
8'h05 : rvCrc[17] <= 32'h8d7ab4cf;
8'h06 : rvCrc[17] <= 32'h0a13d3e7;
8'h07 : rvCrc[17] <= 32'h8b740592;
8'h08 : rvCrc[17] <= 32'h183ac574;
8'h09 : rvCrc[17] <= 32'h995d1301;
8'h0a : rvCrc[17] <= 32'h1e347429;
8'h0b : rvCrc[17] <= 32'h9f53a25c;
8'h0c : rvCrc[17] <= 32'h1427a7ce;
8'h0d : rvCrc[17] <= 32'h954071bb;
8'h0e : rvCrc[17] <= 32'h12291693;
8'h0f : rvCrc[17] <= 32'h934ec0e6;
8'h10 : rvCrc[17] <= 32'h30758ae8;
8'h11 : rvCrc[17] <= 32'hb1125c9d;
8'h12 : rvCrc[17] <= 32'h367b3bb5;
8'h13 : rvCrc[17] <= 32'hb71cedc0;
8'h14 : rvCrc[17] <= 32'h3c68e852;
8'h15 : rvCrc[17] <= 32'hbd0f3e27;
8'h16 : rvCrc[17] <= 32'h3a66590f;
8'h17 : rvCrc[17] <= 32'hbb018f7a;
8'h18 : rvCrc[17] <= 32'h284f4f9c;
8'h19 : rvCrc[17] <= 32'ha92899e9;
8'h1a : rvCrc[17] <= 32'h2e41fec1;
8'h1b : rvCrc[17] <= 32'haf2628b4;
8'h1c : rvCrc[17] <= 32'h24522d26;
8'h1d : rvCrc[17] <= 32'ha535fb53;
8'h1e : rvCrc[17] <= 32'h225c9c7b;
8'h1f : rvCrc[17] <= 32'ha33b4a0e;
8'h20 : rvCrc[17] <= 32'h60eb15d0;
8'h21 : rvCrc[17] <= 32'he18cc3a5;
8'h22 : rvCrc[17] <= 32'h66e5a48d;
8'h23 : rvCrc[17] <= 32'he78272f8;
8'h24 : rvCrc[17] <= 32'h6cf6776a;
8'h25 : rvCrc[17] <= 32'hed91a11f;
8'h26 : rvCrc[17] <= 32'h6af8c637;
8'h27 : rvCrc[17] <= 32'heb9f1042;
8'h28 : rvCrc[17] <= 32'h78d1d0a4;
8'h29 : rvCrc[17] <= 32'hf9b606d1;
8'h2a : rvCrc[17] <= 32'h7edf61f9;
8'h2b : rvCrc[17] <= 32'hffb8b78c;
8'h2c : rvCrc[17] <= 32'h74ccb21e;
8'h2d : rvCrc[17] <= 32'hf5ab646b;
8'h2e : rvCrc[17] <= 32'h72c20343;
8'h2f : rvCrc[17] <= 32'hf3a5d536;
8'h30 : rvCrc[17] <= 32'h509e9f38;
8'h31 : rvCrc[17] <= 32'hd1f9494d;
8'h32 : rvCrc[17] <= 32'h56902e65;
8'h33 : rvCrc[17] <= 32'hd7f7f810;
8'h34 : rvCrc[17] <= 32'h5c83fd82;
8'h35 : rvCrc[17] <= 32'hdde42bf7;
8'h36 : rvCrc[17] <= 32'h5a8d4cdf;
8'h37 : rvCrc[17] <= 32'hdbea9aaa;
8'h38 : rvCrc[17] <= 32'h48a45a4c;
8'h39 : rvCrc[17] <= 32'hc9c38c39;
8'h3a : rvCrc[17] <= 32'h4eaaeb11;
8'h3b : rvCrc[17] <= 32'hcfcd3d64;
8'h3c : rvCrc[17] <= 32'h44b938f6;
8'h3d : rvCrc[17] <= 32'hc5deee83;
8'h3e : rvCrc[17] <= 32'h42b789ab;
8'h3f : rvCrc[17] <= 32'hc3d05fde;
8'h40 : rvCrc[17] <= 32'hc1d62ba0;
8'h41 : rvCrc[17] <= 32'h40b1fdd5;
8'h42 : rvCrc[17] <= 32'hc7d89afd;
8'h43 : rvCrc[17] <= 32'h46bf4c88;
8'h44 : rvCrc[17] <= 32'hcdcb491a;
8'h45 : rvCrc[17] <= 32'h4cac9f6f;
8'h46 : rvCrc[17] <= 32'hcbc5f847;
8'h47 : rvCrc[17] <= 32'h4aa22e32;
8'h48 : rvCrc[17] <= 32'hd9eceed4;
8'h49 : rvCrc[17] <= 32'h588b38a1;
8'h4a : rvCrc[17] <= 32'hdfe25f89;
8'h4b : rvCrc[17] <= 32'h5e8589fc;
8'h4c : rvCrc[17] <= 32'hd5f18c6e;
8'h4d : rvCrc[17] <= 32'h54965a1b;
8'h4e : rvCrc[17] <= 32'hd3ff3d33;
8'h4f : rvCrc[17] <= 32'h5298eb46;
8'h50 : rvCrc[17] <= 32'hf1a3a148;
8'h51 : rvCrc[17] <= 32'h70c4773d;
8'h52 : rvCrc[17] <= 32'hf7ad1015;
8'h53 : rvCrc[17] <= 32'h76cac660;
8'h54 : rvCrc[17] <= 32'hfdbec3f2;
8'h55 : rvCrc[17] <= 32'h7cd91587;
8'h56 : rvCrc[17] <= 32'hfbb072af;
8'h57 : rvCrc[17] <= 32'h7ad7a4da;
8'h58 : rvCrc[17] <= 32'he999643c;
8'h59 : rvCrc[17] <= 32'h68feb249;
8'h5a : rvCrc[17] <= 32'hef97d561;
8'h5b : rvCrc[17] <= 32'h6ef00314;
8'h5c : rvCrc[17] <= 32'he5840686;
8'h5d : rvCrc[17] <= 32'h64e3d0f3;
8'h5e : rvCrc[17] <= 32'he38ab7db;
8'h5f : rvCrc[17] <= 32'h62ed61ae;
8'h60 : rvCrc[17] <= 32'ha13d3e70;
8'h61 : rvCrc[17] <= 32'h205ae805;
8'h62 : rvCrc[17] <= 32'ha7338f2d;
8'h63 : rvCrc[17] <= 32'h26545958;
8'h64 : rvCrc[17] <= 32'had205cca;
8'h65 : rvCrc[17] <= 32'h2c478abf;
8'h66 : rvCrc[17] <= 32'hab2eed97;
8'h67 : rvCrc[17] <= 32'h2a493be2;
8'h68 : rvCrc[17] <= 32'hb907fb04;
8'h69 : rvCrc[17] <= 32'h38602d71;
8'h6a : rvCrc[17] <= 32'hbf094a59;
8'h6b : rvCrc[17] <= 32'h3e6e9c2c;
8'h6c : rvCrc[17] <= 32'hb51a99be;
8'h6d : rvCrc[17] <= 32'h347d4fcb;
8'h6e : rvCrc[17] <= 32'hb31428e3;
8'h6f : rvCrc[17] <= 32'h3273fe96;
8'h70 : rvCrc[17] <= 32'h9148b498;
8'h71 : rvCrc[17] <= 32'h102f62ed;
8'h72 : rvCrc[17] <= 32'h974605c5;
8'h73 : rvCrc[17] <= 32'h1621d3b0;
8'h74 : rvCrc[17] <= 32'h9d55d622;
8'h75 : rvCrc[17] <= 32'h1c320057;
8'h76 : rvCrc[17] <= 32'h9b5b677f;
8'h77 : rvCrc[17] <= 32'h1a3cb10a;
8'h78 : rvCrc[17] <= 32'h897271ec;
8'h79 : rvCrc[17] <= 32'h0815a799;
8'h7a : rvCrc[17] <= 32'h8f7cc0b1;
8'h7b : rvCrc[17] <= 32'h0e1b16c4;
8'h7c : rvCrc[17] <= 32'h856f1356;
8'h7d : rvCrc[17] <= 32'h0408c523;
8'h7e : rvCrc[17] <= 32'h8361a20b;
8'h7f : rvCrc[17] <= 32'h0206747e;
8'h80 : rvCrc[17] <= 32'h876d4af7;
8'h81 : rvCrc[17] <= 32'h060a9c82;
8'h82 : rvCrc[17] <= 32'h8163fbaa;
8'h83 : rvCrc[17] <= 32'h00042ddf;
8'h84 : rvCrc[17] <= 32'h8b70284d;
8'h85 : rvCrc[17] <= 32'h0a17fe38;
8'h86 : rvCrc[17] <= 32'h8d7e9910;
8'h87 : rvCrc[17] <= 32'h0c194f65;
8'h88 : rvCrc[17] <= 32'h9f578f83;
8'h89 : rvCrc[17] <= 32'h1e3059f6;
8'h8a : rvCrc[17] <= 32'h99593ede;
8'h8b : rvCrc[17] <= 32'h183ee8ab;
8'h8c : rvCrc[17] <= 32'h934aed39;
8'h8d : rvCrc[17] <= 32'h122d3b4c;
8'h8e : rvCrc[17] <= 32'h95445c64;
8'h8f : rvCrc[17] <= 32'h14238a11;
8'h90 : rvCrc[17] <= 32'hb718c01f;
8'h91 : rvCrc[17] <= 32'h367f166a;
8'h92 : rvCrc[17] <= 32'hb1167142;
8'h93 : rvCrc[17] <= 32'h3071a737;
8'h94 : rvCrc[17] <= 32'hbb05a2a5;
8'h95 : rvCrc[17] <= 32'h3a6274d0;
8'h96 : rvCrc[17] <= 32'hbd0b13f8;
8'h97 : rvCrc[17] <= 32'h3c6cc58d;
8'h98 : rvCrc[17] <= 32'haf22056b;
8'h99 : rvCrc[17] <= 32'h2e45d31e;
8'h9a : rvCrc[17] <= 32'ha92cb436;
8'h9b : rvCrc[17] <= 32'h284b6243;
8'h9c : rvCrc[17] <= 32'ha33f67d1;
8'h9d : rvCrc[17] <= 32'h2258b1a4;
8'h9e : rvCrc[17] <= 32'ha531d68c;
8'h9f : rvCrc[17] <= 32'h245600f9;
8'ha0 : rvCrc[17] <= 32'he7865f27;
8'ha1 : rvCrc[17] <= 32'h66e18952;
8'ha2 : rvCrc[17] <= 32'he188ee7a;
8'ha3 : rvCrc[17] <= 32'h60ef380f;
8'ha4 : rvCrc[17] <= 32'heb9b3d9d;
8'ha5 : rvCrc[17] <= 32'h6afcebe8;
8'ha6 : rvCrc[17] <= 32'hed958cc0;
8'ha7 : rvCrc[17] <= 32'h6cf25ab5;
8'ha8 : rvCrc[17] <= 32'hffbc9a53;
8'ha9 : rvCrc[17] <= 32'h7edb4c26;
8'haa : rvCrc[17] <= 32'hf9b22b0e;
8'hab : rvCrc[17] <= 32'h78d5fd7b;
8'hac : rvCrc[17] <= 32'hf3a1f8e9;
8'had : rvCrc[17] <= 32'h72c62e9c;
8'hae : rvCrc[17] <= 32'hf5af49b4;
8'haf : rvCrc[17] <= 32'h74c89fc1;
8'hb0 : rvCrc[17] <= 32'hd7f3d5cf;
8'hb1 : rvCrc[17] <= 32'h569403ba;
8'hb2 : rvCrc[17] <= 32'hd1fd6492;
8'hb3 : rvCrc[17] <= 32'h509ab2e7;
8'hb4 : rvCrc[17] <= 32'hdbeeb775;
8'hb5 : rvCrc[17] <= 32'h5a896100;
8'hb6 : rvCrc[17] <= 32'hdde00628;
8'hb7 : rvCrc[17] <= 32'h5c87d05d;
8'hb8 : rvCrc[17] <= 32'hcfc910bb;
8'hb9 : rvCrc[17] <= 32'h4eaec6ce;
8'hba : rvCrc[17] <= 32'hc9c7a1e6;
8'hbb : rvCrc[17] <= 32'h48a07793;
8'hbc : rvCrc[17] <= 32'hc3d47201;
8'hbd : rvCrc[17] <= 32'h42b3a474;
8'hbe : rvCrc[17] <= 32'hc5dac35c;
8'hbf : rvCrc[17] <= 32'h44bd1529;
8'hc0 : rvCrc[17] <= 32'h46bb6157;
8'hc1 : rvCrc[17] <= 32'hc7dcb722;
8'hc2 : rvCrc[17] <= 32'h40b5d00a;
8'hc3 : rvCrc[17] <= 32'hc1d2067f;
8'hc4 : rvCrc[17] <= 32'h4aa603ed;
8'hc5 : rvCrc[17] <= 32'hcbc1d598;
8'hc6 : rvCrc[17] <= 32'h4ca8b2b0;
8'hc7 : rvCrc[17] <= 32'hcdcf64c5;
8'hc8 : rvCrc[17] <= 32'h5e81a423;
8'hc9 : rvCrc[17] <= 32'hdfe67256;
8'hca : rvCrc[17] <= 32'h588f157e;
8'hcb : rvCrc[17] <= 32'hd9e8c30b;
8'hcc : rvCrc[17] <= 32'h529cc699;
8'hcd : rvCrc[17] <= 32'hd3fb10ec;
8'hce : rvCrc[17] <= 32'h549277c4;
8'hcf : rvCrc[17] <= 32'hd5f5a1b1;
8'hd0 : rvCrc[17] <= 32'h76ceebbf;
8'hd1 : rvCrc[17] <= 32'hf7a93dca;
8'hd2 : rvCrc[17] <= 32'h70c05ae2;
8'hd3 : rvCrc[17] <= 32'hf1a78c97;
8'hd4 : rvCrc[17] <= 32'h7ad38905;
8'hd5 : rvCrc[17] <= 32'hfbb45f70;
8'hd6 : rvCrc[17] <= 32'h7cdd3858;
8'hd7 : rvCrc[17] <= 32'hfdbaee2d;
8'hd8 : rvCrc[17] <= 32'h6ef42ecb;
8'hd9 : rvCrc[17] <= 32'hef93f8be;
8'hda : rvCrc[17] <= 32'h68fa9f96;
8'hdb : rvCrc[17] <= 32'he99d49e3;
8'hdc : rvCrc[17] <= 32'h62e94c71;
8'hdd : rvCrc[17] <= 32'he38e9a04;
8'hde : rvCrc[17] <= 32'h64e7fd2c;
8'hdf : rvCrc[17] <= 32'he5802b59;
8'he0 : rvCrc[17] <= 32'h26507487;
8'he1 : rvCrc[17] <= 32'ha737a2f2;
8'he2 : rvCrc[17] <= 32'h205ec5da;
8'he3 : rvCrc[17] <= 32'ha13913af;
8'he4 : rvCrc[17] <= 32'h2a4d163d;
8'he5 : rvCrc[17] <= 32'hab2ac048;
8'he6 : rvCrc[17] <= 32'h2c43a760;
8'he7 : rvCrc[17] <= 32'had247115;
8'he8 : rvCrc[17] <= 32'h3e6ab1f3;
8'he9 : rvCrc[17] <= 32'hbf0d6786;
8'hea : rvCrc[17] <= 32'h386400ae;
8'heb : rvCrc[17] <= 32'hb903d6db;
8'hec : rvCrc[17] <= 32'h3277d349;
8'hed : rvCrc[17] <= 32'hb310053c;
8'hee : rvCrc[17] <= 32'h34796214;
8'hef : rvCrc[17] <= 32'hb51eb461;
8'hf0 : rvCrc[17] <= 32'h1625fe6f;
8'hf1 : rvCrc[17] <= 32'h9742281a;
8'hf2 : rvCrc[17] <= 32'h102b4f32;
8'hf3 : rvCrc[17] <= 32'h914c9947;
8'hf4 : rvCrc[17] <= 32'h1a389cd5;
8'hf5 : rvCrc[17] <= 32'h9b5f4aa0;
8'hf6 : rvCrc[17] <= 32'h1c362d88;
8'hf7 : rvCrc[17] <= 32'h9d51fbfd;
8'hf8 : rvCrc[17] <= 32'h0e1f3b1b;
8'hf9 : rvCrc[17] <= 32'h8f78ed6e;
8'hfa : rvCrc[17] <= 32'h08118a46;
8'hfb : rvCrc[17] <= 32'h89765c33;
8'hfc : rvCrc[17] <= 32'h020259a1;
8'hfd : rvCrc[17] <= 32'h83658fd4;
8'hfe : rvCrc[17] <= 32'h040ce8fc;
8'hff : rvCrc[17] <= 32'h856b3e89;
endcase
case(iv_Input[151:144])
8'h00 : rvCrc[18] <= 32'h00000000;
8'h01 : rvCrc[18] <= 32'h0a1b8859;
8'h02 : rvCrc[18] <= 32'h143710b2;
8'h03 : rvCrc[18] <= 32'h1e2c98eb;
8'h04 : rvCrc[18] <= 32'h286e2164;
8'h05 : rvCrc[18] <= 32'h2275a93d;
8'h06 : rvCrc[18] <= 32'h3c5931d6;
8'h07 : rvCrc[18] <= 32'h3642b98f;
8'h08 : rvCrc[18] <= 32'h50dc42c8;
8'h09 : rvCrc[18] <= 32'h5ac7ca91;
8'h0a : rvCrc[18] <= 32'h44eb527a;
8'h0b : rvCrc[18] <= 32'h4ef0da23;
8'h0c : rvCrc[18] <= 32'h78b263ac;
8'h0d : rvCrc[18] <= 32'h72a9ebf5;
8'h0e : rvCrc[18] <= 32'h6c85731e;
8'h0f : rvCrc[18] <= 32'h669efb47;
8'h10 : rvCrc[18] <= 32'ha1b88590;
8'h11 : rvCrc[18] <= 32'haba30dc9;
8'h12 : rvCrc[18] <= 32'hb58f9522;
8'h13 : rvCrc[18] <= 32'hbf941d7b;
8'h14 : rvCrc[18] <= 32'h89d6a4f4;
8'h15 : rvCrc[18] <= 32'h83cd2cad;
8'h16 : rvCrc[18] <= 32'h9de1b446;
8'h17 : rvCrc[18] <= 32'h97fa3c1f;
8'h18 : rvCrc[18] <= 32'hf164c758;
8'h19 : rvCrc[18] <= 32'hfb7f4f01;
8'h1a : rvCrc[18] <= 32'he553d7ea;
8'h1b : rvCrc[18] <= 32'hef485fb3;
8'h1c : rvCrc[18] <= 32'hd90ae63c;
8'h1d : rvCrc[18] <= 32'hd3116e65;
8'h1e : rvCrc[18] <= 32'hcd3df68e;
8'h1f : rvCrc[18] <= 32'hc7267ed7;
8'h20 : rvCrc[18] <= 32'h47b01697;
8'h21 : rvCrc[18] <= 32'h4dab9ece;
8'h22 : rvCrc[18] <= 32'h53870625;
8'h23 : rvCrc[18] <= 32'h599c8e7c;
8'h24 : rvCrc[18] <= 32'h6fde37f3;
8'h25 : rvCrc[18] <= 32'h65c5bfaa;
8'h26 : rvCrc[18] <= 32'h7be92741;
8'h27 : rvCrc[18] <= 32'h71f2af18;
8'h28 : rvCrc[18] <= 32'h176c545f;
8'h29 : rvCrc[18] <= 32'h1d77dc06;
8'h2a : rvCrc[18] <= 32'h035b44ed;
8'h2b : rvCrc[18] <= 32'h0940ccb4;
8'h2c : rvCrc[18] <= 32'h3f02753b;
8'h2d : rvCrc[18] <= 32'h3519fd62;
8'h2e : rvCrc[18] <= 32'h2b356589;
8'h2f : rvCrc[18] <= 32'h212eedd0;
8'h30 : rvCrc[18] <= 32'he6089307;
8'h31 : rvCrc[18] <= 32'hec131b5e;
8'h32 : rvCrc[18] <= 32'hf23f83b5;
8'h33 : rvCrc[18] <= 32'hf8240bec;
8'h34 : rvCrc[18] <= 32'hce66b263;
8'h35 : rvCrc[18] <= 32'hc47d3a3a;
8'h36 : rvCrc[18] <= 32'hda51a2d1;
8'h37 : rvCrc[18] <= 32'hd04a2a88;
8'h38 : rvCrc[18] <= 32'hb6d4d1cf;
8'h39 : rvCrc[18] <= 32'hbccf5996;
8'h3a : rvCrc[18] <= 32'ha2e3c17d;
8'h3b : rvCrc[18] <= 32'ha8f84924;
8'h3c : rvCrc[18] <= 32'h9ebaf0ab;
8'h3d : rvCrc[18] <= 32'h94a178f2;
8'h3e : rvCrc[18] <= 32'h8a8de019;
8'h3f : rvCrc[18] <= 32'h80966840;
8'h40 : rvCrc[18] <= 32'h8f602d2e;
8'h41 : rvCrc[18] <= 32'h857ba577;
8'h42 : rvCrc[18] <= 32'h9b573d9c;
8'h43 : rvCrc[18] <= 32'h914cb5c5;
8'h44 : rvCrc[18] <= 32'ha70e0c4a;
8'h45 : rvCrc[18] <= 32'had158413;
8'h46 : rvCrc[18] <= 32'hb3391cf8;
8'h47 : rvCrc[18] <= 32'hb92294a1;
8'h48 : rvCrc[18] <= 32'hdfbc6fe6;
8'h49 : rvCrc[18] <= 32'hd5a7e7bf;
8'h4a : rvCrc[18] <= 32'hcb8b7f54;
8'h4b : rvCrc[18] <= 32'hc190f70d;
8'h4c : rvCrc[18] <= 32'hf7d24e82;
8'h4d : rvCrc[18] <= 32'hfdc9c6db;
8'h4e : rvCrc[18] <= 32'he3e55e30;
8'h4f : rvCrc[18] <= 32'he9fed669;
8'h50 : rvCrc[18] <= 32'h2ed8a8be;
8'h51 : rvCrc[18] <= 32'h24c320e7;
8'h52 : rvCrc[18] <= 32'h3aefb80c;
8'h53 : rvCrc[18] <= 32'h30f43055;
8'h54 : rvCrc[18] <= 32'h06b689da;
8'h55 : rvCrc[18] <= 32'h0cad0183;
8'h56 : rvCrc[18] <= 32'h12819968;
8'h57 : rvCrc[18] <= 32'h189a1131;
8'h58 : rvCrc[18] <= 32'h7e04ea76;
8'h59 : rvCrc[18] <= 32'h741f622f;
8'h5a : rvCrc[18] <= 32'h6a33fac4;
8'h5b : rvCrc[18] <= 32'h6028729d;
8'h5c : rvCrc[18] <= 32'h566acb12;
8'h5d : rvCrc[18] <= 32'h5c71434b;
8'h5e : rvCrc[18] <= 32'h425ddba0;
8'h5f : rvCrc[18] <= 32'h484653f9;
8'h60 : rvCrc[18] <= 32'hc8d03bb9;
8'h61 : rvCrc[18] <= 32'hc2cbb3e0;
8'h62 : rvCrc[18] <= 32'hdce72b0b;
8'h63 : rvCrc[18] <= 32'hd6fca352;
8'h64 : rvCrc[18] <= 32'he0be1add;
8'h65 : rvCrc[18] <= 32'heaa59284;
8'h66 : rvCrc[18] <= 32'hf4890a6f;
8'h67 : rvCrc[18] <= 32'hfe928236;
8'h68 : rvCrc[18] <= 32'h980c7971;
8'h69 : rvCrc[18] <= 32'h9217f128;
8'h6a : rvCrc[18] <= 32'h8c3b69c3;
8'h6b : rvCrc[18] <= 32'h8620e19a;
8'h6c : rvCrc[18] <= 32'hb0625815;
8'h6d : rvCrc[18] <= 32'hba79d04c;
8'h6e : rvCrc[18] <= 32'ha45548a7;
8'h6f : rvCrc[18] <= 32'hae4ec0fe;
8'h70 : rvCrc[18] <= 32'h6968be29;
8'h71 : rvCrc[18] <= 32'h63733670;
8'h72 : rvCrc[18] <= 32'h7d5fae9b;
8'h73 : rvCrc[18] <= 32'h774426c2;
8'h74 : rvCrc[18] <= 32'h41069f4d;
8'h75 : rvCrc[18] <= 32'h4b1d1714;
8'h76 : rvCrc[18] <= 32'h55318fff;
8'h77 : rvCrc[18] <= 32'h5f2a07a6;
8'h78 : rvCrc[18] <= 32'h39b4fce1;
8'h79 : rvCrc[18] <= 32'h33af74b8;
8'h7a : rvCrc[18] <= 32'h2d83ec53;
8'h7b : rvCrc[18] <= 32'h2798640a;
8'h7c : rvCrc[18] <= 32'h11dadd85;
8'h7d : rvCrc[18] <= 32'h1bc155dc;
8'h7e : rvCrc[18] <= 32'h05edcd37;
8'h7f : rvCrc[18] <= 32'h0ff6456e;
8'h80 : rvCrc[18] <= 32'h1a0147eb;
8'h81 : rvCrc[18] <= 32'h101acfb2;
8'h82 : rvCrc[18] <= 32'h0e365759;
8'h83 : rvCrc[18] <= 32'h042ddf00;
8'h84 : rvCrc[18] <= 32'h326f668f;
8'h85 : rvCrc[18] <= 32'h3874eed6;
8'h86 : rvCrc[18] <= 32'h2658763d;
8'h87 : rvCrc[18] <= 32'h2c43fe64;
8'h88 : rvCrc[18] <= 32'h4add0523;
8'h89 : rvCrc[18] <= 32'h40c68d7a;
8'h8a : rvCrc[18] <= 32'h5eea1591;
8'h8b : rvCrc[18] <= 32'h54f19dc8;
8'h8c : rvCrc[18] <= 32'h62b32447;
8'h8d : rvCrc[18] <= 32'h68a8ac1e;
8'h8e : rvCrc[18] <= 32'h768434f5;
8'h8f : rvCrc[18] <= 32'h7c9fbcac;
8'h90 : rvCrc[18] <= 32'hbbb9c27b;
8'h91 : rvCrc[18] <= 32'hb1a24a22;
8'h92 : rvCrc[18] <= 32'haf8ed2c9;
8'h93 : rvCrc[18] <= 32'ha5955a90;
8'h94 : rvCrc[18] <= 32'h93d7e31f;
8'h95 : rvCrc[18] <= 32'h99cc6b46;
8'h96 : rvCrc[18] <= 32'h87e0f3ad;
8'h97 : rvCrc[18] <= 32'h8dfb7bf4;
8'h98 : rvCrc[18] <= 32'heb6580b3;
8'h99 : rvCrc[18] <= 32'he17e08ea;
8'h9a : rvCrc[18] <= 32'hff529001;
8'h9b : rvCrc[18] <= 32'hf5491858;
8'h9c : rvCrc[18] <= 32'hc30ba1d7;
8'h9d : rvCrc[18] <= 32'hc910298e;
8'h9e : rvCrc[18] <= 32'hd73cb165;
8'h9f : rvCrc[18] <= 32'hdd27393c;
8'ha0 : rvCrc[18] <= 32'h5db1517c;
8'ha1 : rvCrc[18] <= 32'h57aad925;
8'ha2 : rvCrc[18] <= 32'h498641ce;
8'ha3 : rvCrc[18] <= 32'h439dc997;
8'ha4 : rvCrc[18] <= 32'h75df7018;
8'ha5 : rvCrc[18] <= 32'h7fc4f841;
8'ha6 : rvCrc[18] <= 32'h61e860aa;
8'ha7 : rvCrc[18] <= 32'h6bf3e8f3;
8'ha8 : rvCrc[18] <= 32'h0d6d13b4;
8'ha9 : rvCrc[18] <= 32'h07769bed;
8'haa : rvCrc[18] <= 32'h195a0306;
8'hab : rvCrc[18] <= 32'h13418b5f;
8'hac : rvCrc[18] <= 32'h250332d0;
8'had : rvCrc[18] <= 32'h2f18ba89;
8'hae : rvCrc[18] <= 32'h31342262;
8'haf : rvCrc[18] <= 32'h3b2faa3b;
8'hb0 : rvCrc[18] <= 32'hfc09d4ec;
8'hb1 : rvCrc[18] <= 32'hf6125cb5;
8'hb2 : rvCrc[18] <= 32'he83ec45e;
8'hb3 : rvCrc[18] <= 32'he2254c07;
8'hb4 : rvCrc[18] <= 32'hd467f588;
8'hb5 : rvCrc[18] <= 32'hde7c7dd1;
8'hb6 : rvCrc[18] <= 32'hc050e53a;
8'hb7 : rvCrc[18] <= 32'hca4b6d63;
8'hb8 : rvCrc[18] <= 32'hacd59624;
8'hb9 : rvCrc[18] <= 32'ha6ce1e7d;
8'hba : rvCrc[18] <= 32'hb8e28696;
8'hbb : rvCrc[18] <= 32'hb2f90ecf;
8'hbc : rvCrc[18] <= 32'h84bbb740;
8'hbd : rvCrc[18] <= 32'h8ea03f19;
8'hbe : rvCrc[18] <= 32'h908ca7f2;
8'hbf : rvCrc[18] <= 32'h9a972fab;
8'hc0 : rvCrc[18] <= 32'h95616ac5;
8'hc1 : rvCrc[18] <= 32'h9f7ae29c;
8'hc2 : rvCrc[18] <= 32'h81567a77;
8'hc3 : rvCrc[18] <= 32'h8b4df22e;
8'hc4 : rvCrc[18] <= 32'hbd0f4ba1;
8'hc5 : rvCrc[18] <= 32'hb714c3f8;
8'hc6 : rvCrc[18] <= 32'ha9385b13;
8'hc7 : rvCrc[18] <= 32'ha323d34a;
8'hc8 : rvCrc[18] <= 32'hc5bd280d;
8'hc9 : rvCrc[18] <= 32'hcfa6a054;
8'hca : rvCrc[18] <= 32'hd18a38bf;
8'hcb : rvCrc[18] <= 32'hdb91b0e6;
8'hcc : rvCrc[18] <= 32'hedd30969;
8'hcd : rvCrc[18] <= 32'he7c88130;
8'hce : rvCrc[18] <= 32'hf9e419db;
8'hcf : rvCrc[18] <= 32'hf3ff9182;
8'hd0 : rvCrc[18] <= 32'h34d9ef55;
8'hd1 : rvCrc[18] <= 32'h3ec2670c;
8'hd2 : rvCrc[18] <= 32'h20eeffe7;
8'hd3 : rvCrc[18] <= 32'h2af577be;
8'hd4 : rvCrc[18] <= 32'h1cb7ce31;
8'hd5 : rvCrc[18] <= 32'h16ac4668;
8'hd6 : rvCrc[18] <= 32'h0880de83;
8'hd7 : rvCrc[18] <= 32'h029b56da;
8'hd8 : rvCrc[18] <= 32'h6405ad9d;
8'hd9 : rvCrc[18] <= 32'h6e1e25c4;
8'hda : rvCrc[18] <= 32'h7032bd2f;
8'hdb : rvCrc[18] <= 32'h7a293576;
8'hdc : rvCrc[18] <= 32'h4c6b8cf9;
8'hdd : rvCrc[18] <= 32'h467004a0;
8'hde : rvCrc[18] <= 32'h585c9c4b;
8'hdf : rvCrc[18] <= 32'h52471412;
8'he0 : rvCrc[18] <= 32'hd2d17c52;
8'he1 : rvCrc[18] <= 32'hd8caf40b;
8'he2 : rvCrc[18] <= 32'hc6e66ce0;
8'he3 : rvCrc[18] <= 32'hccfde4b9;
8'he4 : rvCrc[18] <= 32'hfabf5d36;
8'he5 : rvCrc[18] <= 32'hf0a4d56f;
8'he6 : rvCrc[18] <= 32'hee884d84;
8'he7 : rvCrc[18] <= 32'he493c5dd;
8'he8 : rvCrc[18] <= 32'h820d3e9a;
8'he9 : rvCrc[18] <= 32'h8816b6c3;
8'hea : rvCrc[18] <= 32'h963a2e28;
8'heb : rvCrc[18] <= 32'h9c21a671;
8'hec : rvCrc[18] <= 32'haa631ffe;
8'hed : rvCrc[18] <= 32'ha07897a7;
8'hee : rvCrc[18] <= 32'hbe540f4c;
8'hef : rvCrc[18] <= 32'hb44f8715;
8'hf0 : rvCrc[18] <= 32'h7369f9c2;
8'hf1 : rvCrc[18] <= 32'h7972719b;
8'hf2 : rvCrc[18] <= 32'h675ee970;
8'hf3 : rvCrc[18] <= 32'h6d456129;
8'hf4 : rvCrc[18] <= 32'h5b07d8a6;
8'hf5 : rvCrc[18] <= 32'h511c50ff;
8'hf6 : rvCrc[18] <= 32'h4f30c814;
8'hf7 : rvCrc[18] <= 32'h452b404d;
8'hf8 : rvCrc[18] <= 32'h23b5bb0a;
8'hf9 : rvCrc[18] <= 32'h29ae3353;
8'hfa : rvCrc[18] <= 32'h3782abb8;
8'hfb : rvCrc[18] <= 32'h3d9923e1;
8'hfc : rvCrc[18] <= 32'h0bdb9a6e;
8'hfd : rvCrc[18] <= 32'h01c01237;
8'hfe : rvCrc[18] <= 32'h1fec8adc;
8'hff : rvCrc[18] <= 32'h15f70285;
endcase
case(iv_Input[159:152])
8'h00 : rvCrc[19] <= 32'h00000000;
8'h01 : rvCrc[19] <= 32'h34028fd6;
8'h02 : rvCrc[19] <= 32'h68051fac;
8'h03 : rvCrc[19] <= 32'h5c07907a;
8'h04 : rvCrc[19] <= 32'hd00a3f58;
8'h05 : rvCrc[19] <= 32'he408b08e;
8'h06 : rvCrc[19] <= 32'hb80f20f4;
8'h07 : rvCrc[19] <= 32'h8c0daf22;
8'h08 : rvCrc[19] <= 32'ha4d56307;
8'h09 : rvCrc[19] <= 32'h90d7ecd1;
8'h0a : rvCrc[19] <= 32'hccd07cab;
8'h0b : rvCrc[19] <= 32'hf8d2f37d;
8'h0c : rvCrc[19] <= 32'h74df5c5f;
8'h0d : rvCrc[19] <= 32'h40ddd389;
8'h0e : rvCrc[19] <= 32'h1cda43f3;
8'h0f : rvCrc[19] <= 32'h28d8cc25;
8'h10 : rvCrc[19] <= 32'h4d6bdbb9;
8'h11 : rvCrc[19] <= 32'h7969546f;
8'h12 : rvCrc[19] <= 32'h256ec415;
8'h13 : rvCrc[19] <= 32'h116c4bc3;
8'h14 : rvCrc[19] <= 32'h9d61e4e1;
8'h15 : rvCrc[19] <= 32'ha9636b37;
8'h16 : rvCrc[19] <= 32'hf564fb4d;
8'h17 : rvCrc[19] <= 32'hc166749b;
8'h18 : rvCrc[19] <= 32'he9beb8be;
8'h19 : rvCrc[19] <= 32'hddbc3768;
8'h1a : rvCrc[19] <= 32'h81bba712;
8'h1b : rvCrc[19] <= 32'hb5b928c4;
8'h1c : rvCrc[19] <= 32'h39b487e6;
8'h1d : rvCrc[19] <= 32'h0db60830;
8'h1e : rvCrc[19] <= 32'h51b1984a;
8'h1f : rvCrc[19] <= 32'h65b3179c;
8'h20 : rvCrc[19] <= 32'h9ad7b772;
8'h21 : rvCrc[19] <= 32'haed538a4;
8'h22 : rvCrc[19] <= 32'hf2d2a8de;
8'h23 : rvCrc[19] <= 32'hc6d02708;
8'h24 : rvCrc[19] <= 32'h4add882a;
8'h25 : rvCrc[19] <= 32'h7edf07fc;
8'h26 : rvCrc[19] <= 32'h22d89786;
8'h27 : rvCrc[19] <= 32'h16da1850;
8'h28 : rvCrc[19] <= 32'h3e02d475;
8'h29 : rvCrc[19] <= 32'h0a005ba3;
8'h2a : rvCrc[19] <= 32'h5607cbd9;
8'h2b : rvCrc[19] <= 32'h6205440f;
8'h2c : rvCrc[19] <= 32'hee08eb2d;
8'h2d : rvCrc[19] <= 32'hda0a64fb;
8'h2e : rvCrc[19] <= 32'h860df481;
8'h2f : rvCrc[19] <= 32'hb20f7b57;
8'h30 : rvCrc[19] <= 32'hd7bc6ccb;
8'h31 : rvCrc[19] <= 32'he3bee31d;
8'h32 : rvCrc[19] <= 32'hbfb97367;
8'h33 : rvCrc[19] <= 32'h8bbbfcb1;
8'h34 : rvCrc[19] <= 32'h07b65393;
8'h35 : rvCrc[19] <= 32'h33b4dc45;
8'h36 : rvCrc[19] <= 32'h6fb34c3f;
8'h37 : rvCrc[19] <= 32'h5bb1c3e9;
8'h38 : rvCrc[19] <= 32'h73690fcc;
8'h39 : rvCrc[19] <= 32'h476b801a;
8'h3a : rvCrc[19] <= 32'h1b6c1060;
8'h3b : rvCrc[19] <= 32'h2f6e9fb6;
8'h3c : rvCrc[19] <= 32'ha3633094;
8'h3d : rvCrc[19] <= 32'h9761bf42;
8'h3e : rvCrc[19] <= 32'hcb662f38;
8'h3f : rvCrc[19] <= 32'hff64a0ee;
8'h40 : rvCrc[19] <= 32'h316e7353;
8'h41 : rvCrc[19] <= 32'h056cfc85;
8'h42 : rvCrc[19] <= 32'h596b6cff;
8'h43 : rvCrc[19] <= 32'h6d69e329;
8'h44 : rvCrc[19] <= 32'he1644c0b;
8'h45 : rvCrc[19] <= 32'hd566c3dd;
8'h46 : rvCrc[19] <= 32'h896153a7;
8'h47 : rvCrc[19] <= 32'hbd63dc71;
8'h48 : rvCrc[19] <= 32'h95bb1054;
8'h49 : rvCrc[19] <= 32'ha1b99f82;
8'h4a : rvCrc[19] <= 32'hfdbe0ff8;
8'h4b : rvCrc[19] <= 32'hc9bc802e;
8'h4c : rvCrc[19] <= 32'h45b12f0c;
8'h4d : rvCrc[19] <= 32'h71b3a0da;
8'h4e : rvCrc[19] <= 32'h2db430a0;
8'h4f : rvCrc[19] <= 32'h19b6bf76;
8'h50 : rvCrc[19] <= 32'h7c05a8ea;
8'h51 : rvCrc[19] <= 32'h4807273c;
8'h52 : rvCrc[19] <= 32'h1400b746;
8'h53 : rvCrc[19] <= 32'h20023890;
8'h54 : rvCrc[19] <= 32'hac0f97b2;
8'h55 : rvCrc[19] <= 32'h980d1864;
8'h56 : rvCrc[19] <= 32'hc40a881e;
8'h57 : rvCrc[19] <= 32'hf00807c8;
8'h58 : rvCrc[19] <= 32'hd8d0cbed;
8'h59 : rvCrc[19] <= 32'hecd2443b;
8'h5a : rvCrc[19] <= 32'hb0d5d441;
8'h5b : rvCrc[19] <= 32'h84d75b97;
8'h5c : rvCrc[19] <= 32'h08daf4b5;
8'h5d : rvCrc[19] <= 32'h3cd87b63;
8'h5e : rvCrc[19] <= 32'h60dfeb19;
8'h5f : rvCrc[19] <= 32'h54dd64cf;
8'h60 : rvCrc[19] <= 32'habb9c421;
8'h61 : rvCrc[19] <= 32'h9fbb4bf7;
8'h62 : rvCrc[19] <= 32'hc3bcdb8d;
8'h63 : rvCrc[19] <= 32'hf7be545b;
8'h64 : rvCrc[19] <= 32'h7bb3fb79;
8'h65 : rvCrc[19] <= 32'h4fb174af;
8'h66 : rvCrc[19] <= 32'h13b6e4d5;
8'h67 : rvCrc[19] <= 32'h27b46b03;
8'h68 : rvCrc[19] <= 32'h0f6ca726;
8'h69 : rvCrc[19] <= 32'h3b6e28f0;
8'h6a : rvCrc[19] <= 32'h6769b88a;
8'h6b : rvCrc[19] <= 32'h536b375c;
8'h6c : rvCrc[19] <= 32'hdf66987e;
8'h6d : rvCrc[19] <= 32'heb6417a8;
8'h6e : rvCrc[19] <= 32'hb76387d2;
8'h6f : rvCrc[19] <= 32'h83610804;
8'h70 : rvCrc[19] <= 32'he6d21f98;
8'h71 : rvCrc[19] <= 32'hd2d0904e;
8'h72 : rvCrc[19] <= 32'h8ed70034;
8'h73 : rvCrc[19] <= 32'hbad58fe2;
8'h74 : rvCrc[19] <= 32'h36d820c0;
8'h75 : rvCrc[19] <= 32'h02daaf16;
8'h76 : rvCrc[19] <= 32'h5edd3f6c;
8'h77 : rvCrc[19] <= 32'h6adfb0ba;
8'h78 : rvCrc[19] <= 32'h42077c9f;
8'h79 : rvCrc[19] <= 32'h7605f349;
8'h7a : rvCrc[19] <= 32'h2a026333;
8'h7b : rvCrc[19] <= 32'h1e00ece5;
8'h7c : rvCrc[19] <= 32'h920d43c7;
8'h7d : rvCrc[19] <= 32'ha60fcc11;
8'h7e : rvCrc[19] <= 32'hfa085c6b;
8'h7f : rvCrc[19] <= 32'hce0ad3bd;
8'h80 : rvCrc[19] <= 32'h62dce6a6;
8'h81 : rvCrc[19] <= 32'h56de6970;
8'h82 : rvCrc[19] <= 32'h0ad9f90a;
8'h83 : rvCrc[19] <= 32'h3edb76dc;
8'h84 : rvCrc[19] <= 32'hb2d6d9fe;
8'h85 : rvCrc[19] <= 32'h86d45628;
8'h86 : rvCrc[19] <= 32'hdad3c652;
8'h87 : rvCrc[19] <= 32'heed14984;
8'h88 : rvCrc[19] <= 32'hc60985a1;
8'h89 : rvCrc[19] <= 32'hf20b0a77;
8'h8a : rvCrc[19] <= 32'hae0c9a0d;
8'h8b : rvCrc[19] <= 32'h9a0e15db;
8'h8c : rvCrc[19] <= 32'h1603baf9;
8'h8d : rvCrc[19] <= 32'h2201352f;
8'h8e : rvCrc[19] <= 32'h7e06a555;
8'h8f : rvCrc[19] <= 32'h4a042a83;
8'h90 : rvCrc[19] <= 32'h2fb73d1f;
8'h91 : rvCrc[19] <= 32'h1bb5b2c9;
8'h92 : rvCrc[19] <= 32'h47b222b3;
8'h93 : rvCrc[19] <= 32'h73b0ad65;
8'h94 : rvCrc[19] <= 32'hffbd0247;
8'h95 : rvCrc[19] <= 32'hcbbf8d91;
8'h96 : rvCrc[19] <= 32'h97b81deb;
8'h97 : rvCrc[19] <= 32'ha3ba923d;
8'h98 : rvCrc[19] <= 32'h8b625e18;
8'h99 : rvCrc[19] <= 32'hbf60d1ce;
8'h9a : rvCrc[19] <= 32'he36741b4;
8'h9b : rvCrc[19] <= 32'hd765ce62;
8'h9c : rvCrc[19] <= 32'h5b686140;
8'h9d : rvCrc[19] <= 32'h6f6aee96;
8'h9e : rvCrc[19] <= 32'h336d7eec;
8'h9f : rvCrc[19] <= 32'h076ff13a;
8'ha0 : rvCrc[19] <= 32'hf80b51d4;
8'ha1 : rvCrc[19] <= 32'hcc09de02;
8'ha2 : rvCrc[19] <= 32'h900e4e78;
8'ha3 : rvCrc[19] <= 32'ha40cc1ae;
8'ha4 : rvCrc[19] <= 32'h28016e8c;
8'ha5 : rvCrc[19] <= 32'h1c03e15a;
8'ha6 : rvCrc[19] <= 32'h40047120;
8'ha7 : rvCrc[19] <= 32'h7406fef6;
8'ha8 : rvCrc[19] <= 32'h5cde32d3;
8'ha9 : rvCrc[19] <= 32'h68dcbd05;
8'haa : rvCrc[19] <= 32'h34db2d7f;
8'hab : rvCrc[19] <= 32'h00d9a2a9;
8'hac : rvCrc[19] <= 32'h8cd40d8b;
8'had : rvCrc[19] <= 32'hb8d6825d;
8'hae : rvCrc[19] <= 32'he4d11227;
8'haf : rvCrc[19] <= 32'hd0d39df1;
8'hb0 : rvCrc[19] <= 32'hb5608a6d;
8'hb1 : rvCrc[19] <= 32'h816205bb;
8'hb2 : rvCrc[19] <= 32'hdd6595c1;
8'hb3 : rvCrc[19] <= 32'he9671a17;
8'hb4 : rvCrc[19] <= 32'h656ab535;
8'hb5 : rvCrc[19] <= 32'h51683ae3;
8'hb6 : rvCrc[19] <= 32'h0d6faa99;
8'hb7 : rvCrc[19] <= 32'h396d254f;
8'hb8 : rvCrc[19] <= 32'h11b5e96a;
8'hb9 : rvCrc[19] <= 32'h25b766bc;
8'hba : rvCrc[19] <= 32'h79b0f6c6;
8'hbb : rvCrc[19] <= 32'h4db27910;
8'hbc : rvCrc[19] <= 32'hc1bfd632;
8'hbd : rvCrc[19] <= 32'hf5bd59e4;
8'hbe : rvCrc[19] <= 32'ha9bac99e;
8'hbf : rvCrc[19] <= 32'h9db84648;
8'hc0 : rvCrc[19] <= 32'h53b295f5;
8'hc1 : rvCrc[19] <= 32'h67b01a23;
8'hc2 : rvCrc[19] <= 32'h3bb78a59;
8'hc3 : rvCrc[19] <= 32'h0fb5058f;
8'hc4 : rvCrc[19] <= 32'h83b8aaad;
8'hc5 : rvCrc[19] <= 32'hb7ba257b;
8'hc6 : rvCrc[19] <= 32'hebbdb501;
8'hc7 : rvCrc[19] <= 32'hdfbf3ad7;
8'hc8 : rvCrc[19] <= 32'hf767f6f2;
8'hc9 : rvCrc[19] <= 32'hc3657924;
8'hca : rvCrc[19] <= 32'h9f62e95e;
8'hcb : rvCrc[19] <= 32'hab606688;
8'hcc : rvCrc[19] <= 32'h276dc9aa;
8'hcd : rvCrc[19] <= 32'h136f467c;
8'hce : rvCrc[19] <= 32'h4f68d606;
8'hcf : rvCrc[19] <= 32'h7b6a59d0;
8'hd0 : rvCrc[19] <= 32'h1ed94e4c;
8'hd1 : rvCrc[19] <= 32'h2adbc19a;
8'hd2 : rvCrc[19] <= 32'h76dc51e0;
8'hd3 : rvCrc[19] <= 32'h42dede36;
8'hd4 : rvCrc[19] <= 32'hced37114;
8'hd5 : rvCrc[19] <= 32'hfad1fec2;
8'hd6 : rvCrc[19] <= 32'ha6d66eb8;
8'hd7 : rvCrc[19] <= 32'h92d4e16e;
8'hd8 : rvCrc[19] <= 32'hba0c2d4b;
8'hd9 : rvCrc[19] <= 32'h8e0ea29d;
8'hda : rvCrc[19] <= 32'hd20932e7;
8'hdb : rvCrc[19] <= 32'he60bbd31;
8'hdc : rvCrc[19] <= 32'h6a061213;
8'hdd : rvCrc[19] <= 32'h5e049dc5;
8'hde : rvCrc[19] <= 32'h02030dbf;
8'hdf : rvCrc[19] <= 32'h36018269;
8'he0 : rvCrc[19] <= 32'hc9652287;
8'he1 : rvCrc[19] <= 32'hfd67ad51;
8'he2 : rvCrc[19] <= 32'ha1603d2b;
8'he3 : rvCrc[19] <= 32'h9562b2fd;
8'he4 : rvCrc[19] <= 32'h196f1ddf;
8'he5 : rvCrc[19] <= 32'h2d6d9209;
8'he6 : rvCrc[19] <= 32'h716a0273;
8'he7 : rvCrc[19] <= 32'h45688da5;
8'he8 : rvCrc[19] <= 32'h6db04180;
8'he9 : rvCrc[19] <= 32'h59b2ce56;
8'hea : rvCrc[19] <= 32'h05b55e2c;
8'heb : rvCrc[19] <= 32'h31b7d1fa;
8'hec : rvCrc[19] <= 32'hbdba7ed8;
8'hed : rvCrc[19] <= 32'h89b8f10e;
8'hee : rvCrc[19] <= 32'hd5bf6174;
8'hef : rvCrc[19] <= 32'he1bdeea2;
8'hf0 : rvCrc[19] <= 32'h840ef93e;
8'hf1 : rvCrc[19] <= 32'hb00c76e8;
8'hf2 : rvCrc[19] <= 32'hec0be692;
8'hf3 : rvCrc[19] <= 32'hd8096944;
8'hf4 : rvCrc[19] <= 32'h5404c666;
8'hf5 : rvCrc[19] <= 32'h600649b0;
8'hf6 : rvCrc[19] <= 32'h3c01d9ca;
8'hf7 : rvCrc[19] <= 32'h0803561c;
8'hf8 : rvCrc[19] <= 32'h20db9a39;
8'hf9 : rvCrc[19] <= 32'h14d915ef;
8'hfa : rvCrc[19] <= 32'h48de8595;
8'hfb : rvCrc[19] <= 32'h7cdc0a43;
8'hfc : rvCrc[19] <= 32'hf0d1a561;
8'hfd : rvCrc[19] <= 32'hc4d32ab7;
8'hfe : rvCrc[19] <= 32'h98d4bacd;
8'hff : rvCrc[19] <= 32'hacd6351b;
endcase
case(iv_Input[167:160])
8'h00 : rvCrc[20] <= 32'h00000000;
8'h01 : rvCrc[20] <= 32'hc5b9cd4c;
8'h02 : rvCrc[20] <= 32'h8fb2872f;
8'h03 : rvCrc[20] <= 32'h4a0b4a63;
8'h04 : rvCrc[20] <= 32'h1ba413e9;
8'h05 : rvCrc[20] <= 32'hde1ddea5;
8'h06 : rvCrc[20] <= 32'h941694c6;
8'h07 : rvCrc[20] <= 32'h51af598a;
8'h08 : rvCrc[20] <= 32'h374827d2;
8'h09 : rvCrc[20] <= 32'hf2f1ea9e;
8'h0a : rvCrc[20] <= 32'hb8faa0fd;
8'h0b : rvCrc[20] <= 32'h7d436db1;
8'h0c : rvCrc[20] <= 32'h2cec343b;
8'h0d : rvCrc[20] <= 32'he955f977;
8'h0e : rvCrc[20] <= 32'ha35eb314;
8'h0f : rvCrc[20] <= 32'h66e77e58;
8'h10 : rvCrc[20] <= 32'h6e904fa4;
8'h11 : rvCrc[20] <= 32'hab2982e8;
8'h12 : rvCrc[20] <= 32'he122c88b;
8'h13 : rvCrc[20] <= 32'h249b05c7;
8'h14 : rvCrc[20] <= 32'h75345c4d;
8'h15 : rvCrc[20] <= 32'hb08d9101;
8'h16 : rvCrc[20] <= 32'hfa86db62;
8'h17 : rvCrc[20] <= 32'h3f3f162e;
8'h18 : rvCrc[20] <= 32'h59d86876;
8'h19 : rvCrc[20] <= 32'h9c61a53a;
8'h1a : rvCrc[20] <= 32'hd66aef59;
8'h1b : rvCrc[20] <= 32'h13d32215;
8'h1c : rvCrc[20] <= 32'h427c7b9f;
8'h1d : rvCrc[20] <= 32'h87c5b6d3;
8'h1e : rvCrc[20] <= 32'hcdcefcb0;
8'h1f : rvCrc[20] <= 32'h087731fc;
8'h20 : rvCrc[20] <= 32'hdd209f48;
8'h21 : rvCrc[20] <= 32'h18995204;
8'h22 : rvCrc[20] <= 32'h52921867;
8'h23 : rvCrc[20] <= 32'h972bd52b;
8'h24 : rvCrc[20] <= 32'hc6848ca1;
8'h25 : rvCrc[20] <= 32'h033d41ed;
8'h26 : rvCrc[20] <= 32'h49360b8e;
8'h27 : rvCrc[20] <= 32'h8c8fc6c2;
8'h28 : rvCrc[20] <= 32'hea68b89a;
8'h29 : rvCrc[20] <= 32'h2fd175d6;
8'h2a : rvCrc[20] <= 32'h65da3fb5;
8'h2b : rvCrc[20] <= 32'ha063f2f9;
8'h2c : rvCrc[20] <= 32'hf1ccab73;
8'h2d : rvCrc[20] <= 32'h3475663f;
8'h2e : rvCrc[20] <= 32'h7e7e2c5c;
8'h2f : rvCrc[20] <= 32'hbbc7e110;
8'h30 : rvCrc[20] <= 32'hb3b0d0ec;
8'h31 : rvCrc[20] <= 32'h76091da0;
8'h32 : rvCrc[20] <= 32'h3c0257c3;
8'h33 : rvCrc[20] <= 32'hf9bb9a8f;
8'h34 : rvCrc[20] <= 32'ha814c305;
8'h35 : rvCrc[20] <= 32'h6dad0e49;
8'h36 : rvCrc[20] <= 32'h27a6442a;
8'h37 : rvCrc[20] <= 32'he21f8966;
8'h38 : rvCrc[20] <= 32'h84f8f73e;
8'h39 : rvCrc[20] <= 32'h41413a72;
8'h3a : rvCrc[20] <= 32'h0b4a7011;
8'h3b : rvCrc[20] <= 32'hcef3bd5d;
8'h3c : rvCrc[20] <= 32'h9f5ce4d7;
8'h3d : rvCrc[20] <= 32'h5ae5299b;
8'h3e : rvCrc[20] <= 32'h10ee63f8;
8'h3f : rvCrc[20] <= 32'hd557aeb4;
8'h40 : rvCrc[20] <= 32'hbe802327;
8'h41 : rvCrc[20] <= 32'h7b39ee6b;
8'h42 : rvCrc[20] <= 32'h3132a408;
8'h43 : rvCrc[20] <= 32'hf48b6944;
8'h44 : rvCrc[20] <= 32'ha52430ce;
8'h45 : rvCrc[20] <= 32'h609dfd82;
8'h46 : rvCrc[20] <= 32'h2a96b7e1;
8'h47 : rvCrc[20] <= 32'hef2f7aad;
8'h48 : rvCrc[20] <= 32'h89c804f5;
8'h49 : rvCrc[20] <= 32'h4c71c9b9;
8'h4a : rvCrc[20] <= 32'h067a83da;
8'h4b : rvCrc[20] <= 32'hc3c34e96;
8'h4c : rvCrc[20] <= 32'h926c171c;
8'h4d : rvCrc[20] <= 32'h57d5da50;
8'h4e : rvCrc[20] <= 32'h1dde9033;
8'h4f : rvCrc[20] <= 32'hd8675d7f;
8'h50 : rvCrc[20] <= 32'hd0106c83;
8'h51 : rvCrc[20] <= 32'h15a9a1cf;
8'h52 : rvCrc[20] <= 32'h5fa2ebac;
8'h53 : rvCrc[20] <= 32'h9a1b26e0;
8'h54 : rvCrc[20] <= 32'hcbb47f6a;
8'h55 : rvCrc[20] <= 32'h0e0db226;
8'h56 : rvCrc[20] <= 32'h4406f845;
8'h57 : rvCrc[20] <= 32'h81bf3509;
8'h58 : rvCrc[20] <= 32'he7584b51;
8'h59 : rvCrc[20] <= 32'h22e1861d;
8'h5a : rvCrc[20] <= 32'h68eacc7e;
8'h5b : rvCrc[20] <= 32'had530132;
8'h5c : rvCrc[20] <= 32'hfcfc58b8;
8'h5d : rvCrc[20] <= 32'h394595f4;
8'h5e : rvCrc[20] <= 32'h734edf97;
8'h5f : rvCrc[20] <= 32'hb6f712db;
8'h60 : rvCrc[20] <= 32'h63a0bc6f;
8'h61 : rvCrc[20] <= 32'ha6197123;
8'h62 : rvCrc[20] <= 32'hec123b40;
8'h63 : rvCrc[20] <= 32'h29abf60c;
8'h64 : rvCrc[20] <= 32'h7804af86;
8'h65 : rvCrc[20] <= 32'hbdbd62ca;
8'h66 : rvCrc[20] <= 32'hf7b628a9;
8'h67 : rvCrc[20] <= 32'h320fe5e5;
8'h68 : rvCrc[20] <= 32'h54e89bbd;
8'h69 : rvCrc[20] <= 32'h915156f1;
8'h6a : rvCrc[20] <= 32'hdb5a1c92;
8'h6b : rvCrc[20] <= 32'h1ee3d1de;
8'h6c : rvCrc[20] <= 32'h4f4c8854;
8'h6d : rvCrc[20] <= 32'h8af54518;
8'h6e : rvCrc[20] <= 32'hc0fe0f7b;
8'h6f : rvCrc[20] <= 32'h0547c237;
8'h70 : rvCrc[20] <= 32'h0d30f3cb;
8'h71 : rvCrc[20] <= 32'hc8893e87;
8'h72 : rvCrc[20] <= 32'h828274e4;
8'h73 : rvCrc[20] <= 32'h473bb9a8;
8'h74 : rvCrc[20] <= 32'h1694e022;
8'h75 : rvCrc[20] <= 32'hd32d2d6e;
8'h76 : rvCrc[20] <= 32'h9926670d;
8'h77 : rvCrc[20] <= 32'h5c9faa41;
8'h78 : rvCrc[20] <= 32'h3a78d419;
8'h79 : rvCrc[20] <= 32'hffc11955;
8'h7a : rvCrc[20] <= 32'hb5ca5336;
8'h7b : rvCrc[20] <= 32'h70739e7a;
8'h7c : rvCrc[20] <= 32'h21dcc7f0;
8'h7d : rvCrc[20] <= 32'he4650abc;
8'h7e : rvCrc[20] <= 32'hae6e40df;
8'h7f : rvCrc[20] <= 32'h6bd78d93;
8'h80 : rvCrc[20] <= 32'h79c15bf9;
8'h81 : rvCrc[20] <= 32'hbc7896b5;
8'h82 : rvCrc[20] <= 32'hf673dcd6;
8'h83 : rvCrc[20] <= 32'h33ca119a;
8'h84 : rvCrc[20] <= 32'h62654810;
8'h85 : rvCrc[20] <= 32'ha7dc855c;
8'h86 : rvCrc[20] <= 32'hedd7cf3f;
8'h87 : rvCrc[20] <= 32'h286e0273;
8'h88 : rvCrc[20] <= 32'h4e897c2b;
8'h89 : rvCrc[20] <= 32'h8b30b167;
8'h8a : rvCrc[20] <= 32'hc13bfb04;
8'h8b : rvCrc[20] <= 32'h04823648;
8'h8c : rvCrc[20] <= 32'h552d6fc2;
8'h8d : rvCrc[20] <= 32'h9094a28e;
8'h8e : rvCrc[20] <= 32'hda9fe8ed;
8'h8f : rvCrc[20] <= 32'h1f2625a1;
8'h90 : rvCrc[20] <= 32'h1751145d;
8'h91 : rvCrc[20] <= 32'hd2e8d911;
8'h92 : rvCrc[20] <= 32'h98e39372;
8'h93 : rvCrc[20] <= 32'h5d5a5e3e;
8'h94 : rvCrc[20] <= 32'h0cf507b4;
8'h95 : rvCrc[20] <= 32'hc94ccaf8;
8'h96 : rvCrc[20] <= 32'h8347809b;
8'h97 : rvCrc[20] <= 32'h46fe4dd7;
8'h98 : rvCrc[20] <= 32'h2019338f;
8'h99 : rvCrc[20] <= 32'he5a0fec3;
8'h9a : rvCrc[20] <= 32'hafabb4a0;
8'h9b : rvCrc[20] <= 32'h6a1279ec;
8'h9c : rvCrc[20] <= 32'h3bbd2066;
8'h9d : rvCrc[20] <= 32'hfe04ed2a;
8'h9e : rvCrc[20] <= 32'hb40fa749;
8'h9f : rvCrc[20] <= 32'h71b66a05;
8'ha0 : rvCrc[20] <= 32'ha4e1c4b1;
8'ha1 : rvCrc[20] <= 32'h615809fd;
8'ha2 : rvCrc[20] <= 32'h2b53439e;
8'ha3 : rvCrc[20] <= 32'heeea8ed2;
8'ha4 : rvCrc[20] <= 32'hbf45d758;
8'ha5 : rvCrc[20] <= 32'h7afc1a14;
8'ha6 : rvCrc[20] <= 32'h30f75077;
8'ha7 : rvCrc[20] <= 32'hf54e9d3b;
8'ha8 : rvCrc[20] <= 32'h93a9e363;
8'ha9 : rvCrc[20] <= 32'h56102e2f;
8'haa : rvCrc[20] <= 32'h1c1b644c;
8'hab : rvCrc[20] <= 32'hd9a2a900;
8'hac : rvCrc[20] <= 32'h880df08a;
8'had : rvCrc[20] <= 32'h4db43dc6;
8'hae : rvCrc[20] <= 32'h07bf77a5;
8'haf : rvCrc[20] <= 32'hc206bae9;
8'hb0 : rvCrc[20] <= 32'hca718b15;
8'hb1 : rvCrc[20] <= 32'h0fc84659;
8'hb2 : rvCrc[20] <= 32'h45c30c3a;
8'hb3 : rvCrc[20] <= 32'h807ac176;
8'hb4 : rvCrc[20] <= 32'hd1d598fc;
8'hb5 : rvCrc[20] <= 32'h146c55b0;
8'hb6 : rvCrc[20] <= 32'h5e671fd3;
8'hb7 : rvCrc[20] <= 32'h9bded29f;
8'hb8 : rvCrc[20] <= 32'hfd39acc7;
8'hb9 : rvCrc[20] <= 32'h3880618b;
8'hba : rvCrc[20] <= 32'h728b2be8;
8'hbb : rvCrc[20] <= 32'hb732e6a4;
8'hbc : rvCrc[20] <= 32'he69dbf2e;
8'hbd : rvCrc[20] <= 32'h23247262;
8'hbe : rvCrc[20] <= 32'h692f3801;
8'hbf : rvCrc[20] <= 32'hac96f54d;
8'hc0 : rvCrc[20] <= 32'hc74178de;
8'hc1 : rvCrc[20] <= 32'h02f8b592;
8'hc2 : rvCrc[20] <= 32'h48f3fff1;
8'hc3 : rvCrc[20] <= 32'h8d4a32bd;
8'hc4 : rvCrc[20] <= 32'hdce56b37;
8'hc5 : rvCrc[20] <= 32'h195ca67b;
8'hc6 : rvCrc[20] <= 32'h5357ec18;
8'hc7 : rvCrc[20] <= 32'h96ee2154;
8'hc8 : rvCrc[20] <= 32'hf0095f0c;
8'hc9 : rvCrc[20] <= 32'h35b09240;
8'hca : rvCrc[20] <= 32'h7fbbd823;
8'hcb : rvCrc[20] <= 32'hba02156f;
8'hcc : rvCrc[20] <= 32'hebad4ce5;
8'hcd : rvCrc[20] <= 32'h2e1481a9;
8'hce : rvCrc[20] <= 32'h641fcbca;
8'hcf : rvCrc[20] <= 32'ha1a60686;
8'hd0 : rvCrc[20] <= 32'ha9d1377a;
8'hd1 : rvCrc[20] <= 32'h6c68fa36;
8'hd2 : rvCrc[20] <= 32'h2663b055;
8'hd3 : rvCrc[20] <= 32'he3da7d19;
8'hd4 : rvCrc[20] <= 32'hb2752493;
8'hd5 : rvCrc[20] <= 32'h77cce9df;
8'hd6 : rvCrc[20] <= 32'h3dc7a3bc;
8'hd7 : rvCrc[20] <= 32'hf87e6ef0;
8'hd8 : rvCrc[20] <= 32'h9e9910a8;
8'hd9 : rvCrc[20] <= 32'h5b20dde4;
8'hda : rvCrc[20] <= 32'h112b9787;
8'hdb : rvCrc[20] <= 32'hd4925acb;
8'hdc : rvCrc[20] <= 32'h853d0341;
8'hdd : rvCrc[20] <= 32'h4084ce0d;
8'hde : rvCrc[20] <= 32'h0a8f846e;
8'hdf : rvCrc[20] <= 32'hcf364922;
8'he0 : rvCrc[20] <= 32'h1a61e796;
8'he1 : rvCrc[20] <= 32'hdfd82ada;
8'he2 : rvCrc[20] <= 32'h95d360b9;
8'he3 : rvCrc[20] <= 32'h506aadf5;
8'he4 : rvCrc[20] <= 32'h01c5f47f;
8'he5 : rvCrc[20] <= 32'hc47c3933;
8'he6 : rvCrc[20] <= 32'h8e777350;
8'he7 : rvCrc[20] <= 32'h4bcebe1c;
8'he8 : rvCrc[20] <= 32'h2d29c044;
8'he9 : rvCrc[20] <= 32'he8900d08;
8'hea : rvCrc[20] <= 32'ha29b476b;
8'heb : rvCrc[20] <= 32'h67228a27;
8'hec : rvCrc[20] <= 32'h368dd3ad;
8'hed : rvCrc[20] <= 32'hf3341ee1;
8'hee : rvCrc[20] <= 32'hb93f5482;
8'hef : rvCrc[20] <= 32'h7c8699ce;
8'hf0 : rvCrc[20] <= 32'h74f1a832;
8'hf1 : rvCrc[20] <= 32'hb148657e;
8'hf2 : rvCrc[20] <= 32'hfb432f1d;
8'hf3 : rvCrc[20] <= 32'h3efae251;
8'hf4 : rvCrc[20] <= 32'h6f55bbdb;
8'hf5 : rvCrc[20] <= 32'haaec7697;
8'hf6 : rvCrc[20] <= 32'he0e73cf4;
8'hf7 : rvCrc[20] <= 32'h255ef1b8;
8'hf8 : rvCrc[20] <= 32'h43b98fe0;
8'hf9 : rvCrc[20] <= 32'h860042ac;
8'hfa : rvCrc[20] <= 32'hcc0b08cf;
8'hfb : rvCrc[20] <= 32'h09b2c583;
8'hfc : rvCrc[20] <= 32'h581d9c09;
8'hfd : rvCrc[20] <= 32'h9da45145;
8'hfe : rvCrc[20] <= 32'hd7af1b26;
8'hff : rvCrc[20] <= 32'h1216d66a;
endcase
case(iv_Input[175:168])
8'h00 : rvCrc[21] <= 32'h00000000;
8'h01 : rvCrc[21] <= 32'hf382b7f2;
8'h02 : rvCrc[21] <= 32'he3c47253;
8'h03 : rvCrc[21] <= 32'h1046c5a1;
8'h04 : rvCrc[21] <= 32'hc349f911;
8'h05 : rvCrc[21] <= 32'h30cb4ee3;
8'h06 : rvCrc[21] <= 32'h208d8b42;
8'h07 : rvCrc[21] <= 32'hd30f3cb0;
8'h08 : rvCrc[21] <= 32'h8252ef95;
8'h09 : rvCrc[21] <= 32'h71d05867;
8'h0a : rvCrc[21] <= 32'h61969dc6;
8'h0b : rvCrc[21] <= 32'h92142a34;
8'h0c : rvCrc[21] <= 32'h411b1684;
8'h0d : rvCrc[21] <= 32'hb299a176;
8'h0e : rvCrc[21] <= 32'ha2df64d7;
8'h0f : rvCrc[21] <= 32'h515dd325;
8'h10 : rvCrc[21] <= 32'h0064c29d;
8'h11 : rvCrc[21] <= 32'hf3e6756f;
8'h12 : rvCrc[21] <= 32'he3a0b0ce;
8'h13 : rvCrc[21] <= 32'h1022073c;
8'h14 : rvCrc[21] <= 32'hc32d3b8c;
8'h15 : rvCrc[21] <= 32'h30af8c7e;
8'h16 : rvCrc[21] <= 32'h20e949df;
8'h17 : rvCrc[21] <= 32'hd36bfe2d;
8'h18 : rvCrc[21] <= 32'h82362d08;
8'h19 : rvCrc[21] <= 32'h71b49afa;
8'h1a : rvCrc[21] <= 32'h61f25f5b;
8'h1b : rvCrc[21] <= 32'h9270e8a9;
8'h1c : rvCrc[21] <= 32'h417fd419;
8'h1d : rvCrc[21] <= 32'hb2fd63eb;
8'h1e : rvCrc[21] <= 32'ha2bba64a;
8'h1f : rvCrc[21] <= 32'h513911b8;
8'h20 : rvCrc[21] <= 32'h00c9853a;
8'h21 : rvCrc[21] <= 32'hf34b32c8;
8'h22 : rvCrc[21] <= 32'he30df769;
8'h23 : rvCrc[21] <= 32'h108f409b;
8'h24 : rvCrc[21] <= 32'hc3807c2b;
8'h25 : rvCrc[21] <= 32'h3002cbd9;
8'h26 : rvCrc[21] <= 32'h20440e78;
8'h27 : rvCrc[21] <= 32'hd3c6b98a;
8'h28 : rvCrc[21] <= 32'h829b6aaf;
8'h29 : rvCrc[21] <= 32'h7119dd5d;
8'h2a : rvCrc[21] <= 32'h615f18fc;
8'h2b : rvCrc[21] <= 32'h92ddaf0e;
8'h2c : rvCrc[21] <= 32'h41d293be;
8'h2d : rvCrc[21] <= 32'hb250244c;
8'h2e : rvCrc[21] <= 32'ha216e1ed;
8'h2f : rvCrc[21] <= 32'h5194561f;
8'h30 : rvCrc[21] <= 32'h00ad47a7;
8'h31 : rvCrc[21] <= 32'hf32ff055;
8'h32 : rvCrc[21] <= 32'he36935f4;
8'h33 : rvCrc[21] <= 32'h10eb8206;
8'h34 : rvCrc[21] <= 32'hc3e4beb6;
8'h35 : rvCrc[21] <= 32'h30660944;
8'h36 : rvCrc[21] <= 32'h2020cce5;
8'h37 : rvCrc[21] <= 32'hd3a27b17;
8'h38 : rvCrc[21] <= 32'h82ffa832;
8'h39 : rvCrc[21] <= 32'h717d1fc0;
8'h3a : rvCrc[21] <= 32'h613bda61;
8'h3b : rvCrc[21] <= 32'h92b96d93;
8'h3c : rvCrc[21] <= 32'h41b65123;
8'h3d : rvCrc[21] <= 32'hb234e6d1;
8'h3e : rvCrc[21] <= 32'ha2722370;
8'h3f : rvCrc[21] <= 32'h51f09482;
8'h40 : rvCrc[21] <= 32'h01930a74;
8'h41 : rvCrc[21] <= 32'hf211bd86;
8'h42 : rvCrc[21] <= 32'he2577827;
8'h43 : rvCrc[21] <= 32'h11d5cfd5;
8'h44 : rvCrc[21] <= 32'hc2daf365;
8'h45 : rvCrc[21] <= 32'h31584497;
8'h46 : rvCrc[21] <= 32'h211e8136;
8'h47 : rvCrc[21] <= 32'hd29c36c4;
8'h48 : rvCrc[21] <= 32'h83c1e5e1;
8'h49 : rvCrc[21] <= 32'h70435213;
8'h4a : rvCrc[21] <= 32'h600597b2;
8'h4b : rvCrc[21] <= 32'h93872040;
8'h4c : rvCrc[21] <= 32'h40881cf0;
8'h4d : rvCrc[21] <= 32'hb30aab02;
8'h4e : rvCrc[21] <= 32'ha34c6ea3;
8'h4f : rvCrc[21] <= 32'h50ced951;
8'h50 : rvCrc[21] <= 32'h01f7c8e9;
8'h51 : rvCrc[21] <= 32'hf2757f1b;
8'h52 : rvCrc[21] <= 32'he233baba;
8'h53 : rvCrc[21] <= 32'h11b10d48;
8'h54 : rvCrc[21] <= 32'hc2be31f8;
8'h55 : rvCrc[21] <= 32'h313c860a;
8'h56 : rvCrc[21] <= 32'h217a43ab;
8'h57 : rvCrc[21] <= 32'hd2f8f459;
8'h58 : rvCrc[21] <= 32'h83a5277c;
8'h59 : rvCrc[21] <= 32'h7027908e;
8'h5a : rvCrc[21] <= 32'h6061552f;
8'h5b : rvCrc[21] <= 32'h93e3e2dd;
8'h5c : rvCrc[21] <= 32'h40ecde6d;
8'h5d : rvCrc[21] <= 32'hb36e699f;
8'h5e : rvCrc[21] <= 32'ha328ac3e;
8'h5f : rvCrc[21] <= 32'h50aa1bcc;
8'h60 : rvCrc[21] <= 32'h015a8f4e;
8'h61 : rvCrc[21] <= 32'hf2d838bc;
8'h62 : rvCrc[21] <= 32'he29efd1d;
8'h63 : rvCrc[21] <= 32'h111c4aef;
8'h64 : rvCrc[21] <= 32'hc213765f;
8'h65 : rvCrc[21] <= 32'h3191c1ad;
8'h66 : rvCrc[21] <= 32'h21d7040c;
8'h67 : rvCrc[21] <= 32'hd255b3fe;
8'h68 : rvCrc[21] <= 32'h830860db;
8'h69 : rvCrc[21] <= 32'h708ad729;
8'h6a : rvCrc[21] <= 32'h60cc1288;
8'h6b : rvCrc[21] <= 32'h934ea57a;
8'h6c : rvCrc[21] <= 32'h404199ca;
8'h6d : rvCrc[21] <= 32'hb3c32e38;
8'h6e : rvCrc[21] <= 32'ha385eb99;
8'h6f : rvCrc[21] <= 32'h50075c6b;
8'h70 : rvCrc[21] <= 32'h013e4dd3;
8'h71 : rvCrc[21] <= 32'hf2bcfa21;
8'h72 : rvCrc[21] <= 32'he2fa3f80;
8'h73 : rvCrc[21] <= 32'h11788872;
8'h74 : rvCrc[21] <= 32'hc277b4c2;
8'h75 : rvCrc[21] <= 32'h31f50330;
8'h76 : rvCrc[21] <= 32'h21b3c691;
8'h77 : rvCrc[21] <= 32'hd2317163;
8'h78 : rvCrc[21] <= 32'h836ca246;
8'h79 : rvCrc[21] <= 32'h70ee15b4;
8'h7a : rvCrc[21] <= 32'h60a8d015;
8'h7b : rvCrc[21] <= 32'h932a67e7;
8'h7c : rvCrc[21] <= 32'h40255b57;
8'h7d : rvCrc[21] <= 32'hb3a7eca5;
8'h7e : rvCrc[21] <= 32'ha3e12904;
8'h7f : rvCrc[21] <= 32'h50639ef6;
8'h80 : rvCrc[21] <= 32'h032614e8;
8'h81 : rvCrc[21] <= 32'hf0a4a31a;
8'h82 : rvCrc[21] <= 32'he0e266bb;
8'h83 : rvCrc[21] <= 32'h1360d149;
8'h84 : rvCrc[21] <= 32'hc06fedf9;
8'h85 : rvCrc[21] <= 32'h33ed5a0b;
8'h86 : rvCrc[21] <= 32'h23ab9faa;
8'h87 : rvCrc[21] <= 32'hd0292858;
8'h88 : rvCrc[21] <= 32'h8174fb7d;
8'h89 : rvCrc[21] <= 32'h72f64c8f;
8'h8a : rvCrc[21] <= 32'h62b0892e;
8'h8b : rvCrc[21] <= 32'h91323edc;
8'h8c : rvCrc[21] <= 32'h423d026c;
8'h8d : rvCrc[21] <= 32'hb1bfb59e;
8'h8e : rvCrc[21] <= 32'ha1f9703f;
8'h8f : rvCrc[21] <= 32'h527bc7cd;
8'h90 : rvCrc[21] <= 32'h0342d675;
8'h91 : rvCrc[21] <= 32'hf0c06187;
8'h92 : rvCrc[21] <= 32'he086a426;
8'h93 : rvCrc[21] <= 32'h130413d4;
8'h94 : rvCrc[21] <= 32'hc00b2f64;
8'h95 : rvCrc[21] <= 32'h33899896;
8'h96 : rvCrc[21] <= 32'h23cf5d37;
8'h97 : rvCrc[21] <= 32'hd04deac5;
8'h98 : rvCrc[21] <= 32'h811039e0;
8'h99 : rvCrc[21] <= 32'h72928e12;
8'h9a : rvCrc[21] <= 32'h62d44bb3;
8'h9b : rvCrc[21] <= 32'h9156fc41;
8'h9c : rvCrc[21] <= 32'h4259c0f1;
8'h9d : rvCrc[21] <= 32'hb1db7703;
8'h9e : rvCrc[21] <= 32'ha19db2a2;
8'h9f : rvCrc[21] <= 32'h521f0550;
8'ha0 : rvCrc[21] <= 32'h03ef91d2;
8'ha1 : rvCrc[21] <= 32'hf06d2620;
8'ha2 : rvCrc[21] <= 32'he02be381;
8'ha3 : rvCrc[21] <= 32'h13a95473;
8'ha4 : rvCrc[21] <= 32'hc0a668c3;
8'ha5 : rvCrc[21] <= 32'h3324df31;
8'ha6 : rvCrc[21] <= 32'h23621a90;
8'ha7 : rvCrc[21] <= 32'hd0e0ad62;
8'ha8 : rvCrc[21] <= 32'h81bd7e47;
8'ha9 : rvCrc[21] <= 32'h723fc9b5;
8'haa : rvCrc[21] <= 32'h62790c14;
8'hab : rvCrc[21] <= 32'h91fbbbe6;
8'hac : rvCrc[21] <= 32'h42f48756;
8'had : rvCrc[21] <= 32'hb17630a4;
8'hae : rvCrc[21] <= 32'ha130f505;
8'haf : rvCrc[21] <= 32'h52b242f7;
8'hb0 : rvCrc[21] <= 32'h038b534f;
8'hb1 : rvCrc[21] <= 32'hf009e4bd;
8'hb2 : rvCrc[21] <= 32'he04f211c;
8'hb3 : rvCrc[21] <= 32'h13cd96ee;
8'hb4 : rvCrc[21] <= 32'hc0c2aa5e;
8'hb5 : rvCrc[21] <= 32'h33401dac;
8'hb6 : rvCrc[21] <= 32'h2306d80d;
8'hb7 : rvCrc[21] <= 32'hd0846fff;
8'hb8 : rvCrc[21] <= 32'h81d9bcda;
8'hb9 : rvCrc[21] <= 32'h725b0b28;
8'hba : rvCrc[21] <= 32'h621dce89;
8'hbb : rvCrc[21] <= 32'h919f797b;
8'hbc : rvCrc[21] <= 32'h429045cb;
8'hbd : rvCrc[21] <= 32'hb112f239;
8'hbe : rvCrc[21] <= 32'ha1543798;
8'hbf : rvCrc[21] <= 32'h52d6806a;
8'hc0 : rvCrc[21] <= 32'h02b51e9c;
8'hc1 : rvCrc[21] <= 32'hf137a96e;
8'hc2 : rvCrc[21] <= 32'he1716ccf;
8'hc3 : rvCrc[21] <= 32'h12f3db3d;
8'hc4 : rvCrc[21] <= 32'hc1fce78d;
8'hc5 : rvCrc[21] <= 32'h327e507f;
8'hc6 : rvCrc[21] <= 32'h223895de;
8'hc7 : rvCrc[21] <= 32'hd1ba222c;
8'hc8 : rvCrc[21] <= 32'h80e7f109;
8'hc9 : rvCrc[21] <= 32'h736546fb;
8'hca : rvCrc[21] <= 32'h6323835a;
8'hcb : rvCrc[21] <= 32'h90a134a8;
8'hcc : rvCrc[21] <= 32'h43ae0818;
8'hcd : rvCrc[21] <= 32'hb02cbfea;
8'hce : rvCrc[21] <= 32'ha06a7a4b;
8'hcf : rvCrc[21] <= 32'h53e8cdb9;
8'hd0 : rvCrc[21] <= 32'h02d1dc01;
8'hd1 : rvCrc[21] <= 32'hf1536bf3;
8'hd2 : rvCrc[21] <= 32'he115ae52;
8'hd3 : rvCrc[21] <= 32'h129719a0;
8'hd4 : rvCrc[21] <= 32'hc1982510;
8'hd5 : rvCrc[21] <= 32'h321a92e2;
8'hd6 : rvCrc[21] <= 32'h225c5743;
8'hd7 : rvCrc[21] <= 32'hd1dee0b1;
8'hd8 : rvCrc[21] <= 32'h80833394;
8'hd9 : rvCrc[21] <= 32'h73018466;
8'hda : rvCrc[21] <= 32'h634741c7;
8'hdb : rvCrc[21] <= 32'h90c5f635;
8'hdc : rvCrc[21] <= 32'h43caca85;
8'hdd : rvCrc[21] <= 32'hb0487d77;
8'hde : rvCrc[21] <= 32'ha00eb8d6;
8'hdf : rvCrc[21] <= 32'h538c0f24;
8'he0 : rvCrc[21] <= 32'h027c9ba6;
8'he1 : rvCrc[21] <= 32'hf1fe2c54;
8'he2 : rvCrc[21] <= 32'he1b8e9f5;
8'he3 : rvCrc[21] <= 32'h123a5e07;
8'he4 : rvCrc[21] <= 32'hc13562b7;
8'he5 : rvCrc[21] <= 32'h32b7d545;
8'he6 : rvCrc[21] <= 32'h22f110e4;
8'he7 : rvCrc[21] <= 32'hd173a716;
8'he8 : rvCrc[21] <= 32'h802e7433;
8'he9 : rvCrc[21] <= 32'h73acc3c1;
8'hea : rvCrc[21] <= 32'h63ea0660;
8'heb : rvCrc[21] <= 32'h9068b192;
8'hec : rvCrc[21] <= 32'h43678d22;
8'hed : rvCrc[21] <= 32'hb0e53ad0;
8'hee : rvCrc[21] <= 32'ha0a3ff71;
8'hef : rvCrc[21] <= 32'h53214883;
8'hf0 : rvCrc[21] <= 32'h0218593b;
8'hf1 : rvCrc[21] <= 32'hf19aeec9;
8'hf2 : rvCrc[21] <= 32'he1dc2b68;
8'hf3 : rvCrc[21] <= 32'h125e9c9a;
8'hf4 : rvCrc[21] <= 32'hc151a02a;
8'hf5 : rvCrc[21] <= 32'h32d317d8;
8'hf6 : rvCrc[21] <= 32'h2295d279;
8'hf7 : rvCrc[21] <= 32'hd117658b;
8'hf8 : rvCrc[21] <= 32'h804ab6ae;
8'hf9 : rvCrc[21] <= 32'h73c8015c;
8'hfa : rvCrc[21] <= 32'h638ec4fd;
8'hfb : rvCrc[21] <= 32'h900c730f;
8'hfc : rvCrc[21] <= 32'h43034fbf;
8'hfd : rvCrc[21] <= 32'hb081f84d;
8'hfe : rvCrc[21] <= 32'ha0c73dec;
8'hff : rvCrc[21] <= 32'h53458a1e;
endcase
case(iv_Input[183:176])
8'h00 : rvCrc[22] <= 32'h00000000;
8'h01 : rvCrc[22] <= 32'h064c29d0;
8'h02 : rvCrc[22] <= 32'h0c9853a0;
8'h03 : rvCrc[22] <= 32'h0ad47a70;
8'h04 : rvCrc[22] <= 32'h1930a740;
8'h05 : rvCrc[22] <= 32'h1f7c8e90;
8'h06 : rvCrc[22] <= 32'h15a8f4e0;
8'h07 : rvCrc[22] <= 32'h13e4dd30;
8'h08 : rvCrc[22] <= 32'h32614e80;
8'h09 : rvCrc[22] <= 32'h342d6750;
8'h0a : rvCrc[22] <= 32'h3ef91d20;
8'h0b : rvCrc[22] <= 32'h38b534f0;
8'h0c : rvCrc[22] <= 32'h2b51e9c0;
8'h0d : rvCrc[22] <= 32'h2d1dc010;
8'h0e : rvCrc[22] <= 32'h27c9ba60;
8'h0f : rvCrc[22] <= 32'h218593b0;
8'h10 : rvCrc[22] <= 32'h64c29d00;
8'h11 : rvCrc[22] <= 32'h628eb4d0;
8'h12 : rvCrc[22] <= 32'h685acea0;
8'h13 : rvCrc[22] <= 32'h6e16e770;
8'h14 : rvCrc[22] <= 32'h7df23a40;
8'h15 : rvCrc[22] <= 32'h7bbe1390;
8'h16 : rvCrc[22] <= 32'h716a69e0;
8'h17 : rvCrc[22] <= 32'h77264030;
8'h18 : rvCrc[22] <= 32'h56a3d380;
8'h19 : rvCrc[22] <= 32'h50effa50;
8'h1a : rvCrc[22] <= 32'h5a3b8020;
8'h1b : rvCrc[22] <= 32'h5c77a9f0;
8'h1c : rvCrc[22] <= 32'h4f9374c0;
8'h1d : rvCrc[22] <= 32'h49df5d10;
8'h1e : rvCrc[22] <= 32'h430b2760;
8'h1f : rvCrc[22] <= 32'h45470eb0;
8'h20 : rvCrc[22] <= 32'hc9853a00;
8'h21 : rvCrc[22] <= 32'hcfc913d0;
8'h22 : rvCrc[22] <= 32'hc51d69a0;
8'h23 : rvCrc[22] <= 32'hc3514070;
8'h24 : rvCrc[22] <= 32'hd0b59d40;
8'h25 : rvCrc[22] <= 32'hd6f9b490;
8'h26 : rvCrc[22] <= 32'hdc2dcee0;
8'h27 : rvCrc[22] <= 32'hda61e730;
8'h28 : rvCrc[22] <= 32'hfbe47480;
8'h29 : rvCrc[22] <= 32'hfda85d50;
8'h2a : rvCrc[22] <= 32'hf77c2720;
8'h2b : rvCrc[22] <= 32'hf1300ef0;
8'h2c : rvCrc[22] <= 32'he2d4d3c0;
8'h2d : rvCrc[22] <= 32'he498fa10;
8'h2e : rvCrc[22] <= 32'hee4c8060;
8'h2f : rvCrc[22] <= 32'he800a9b0;
8'h30 : rvCrc[22] <= 32'had47a700;
8'h31 : rvCrc[22] <= 32'hab0b8ed0;
8'h32 : rvCrc[22] <= 32'ha1dff4a0;
8'h33 : rvCrc[22] <= 32'ha793dd70;
8'h34 : rvCrc[22] <= 32'hb4770040;
8'h35 : rvCrc[22] <= 32'hb23b2990;
8'h36 : rvCrc[22] <= 32'hb8ef53e0;
8'h37 : rvCrc[22] <= 32'hbea37a30;
8'h38 : rvCrc[22] <= 32'h9f26e980;
8'h39 : rvCrc[22] <= 32'h996ac050;
8'h3a : rvCrc[22] <= 32'h93beba20;
8'h3b : rvCrc[22] <= 32'h95f293f0;
8'h3c : rvCrc[22] <= 32'h86164ec0;
8'h3d : rvCrc[22] <= 32'h805a6710;
8'h3e : rvCrc[22] <= 32'h8a8e1d60;
8'h3f : rvCrc[22] <= 32'h8cc234b0;
8'h40 : rvCrc[22] <= 32'h97cb69b7;
8'h41 : rvCrc[22] <= 32'h91874067;
8'h42 : rvCrc[22] <= 32'h9b533a17;
8'h43 : rvCrc[22] <= 32'h9d1f13c7;
8'h44 : rvCrc[22] <= 32'h8efbcef7;
8'h45 : rvCrc[22] <= 32'h88b7e727;
8'h46 : rvCrc[22] <= 32'h82639d57;
8'h47 : rvCrc[22] <= 32'h842fb487;
8'h48 : rvCrc[22] <= 32'ha5aa2737;
8'h49 : rvCrc[22] <= 32'ha3e60ee7;
8'h4a : rvCrc[22] <= 32'ha9327497;
8'h4b : rvCrc[22] <= 32'haf7e5d47;
8'h4c : rvCrc[22] <= 32'hbc9a8077;
8'h4d : rvCrc[22] <= 32'hbad6a9a7;
8'h4e : rvCrc[22] <= 32'hb002d3d7;
8'h4f : rvCrc[22] <= 32'hb64efa07;
8'h50 : rvCrc[22] <= 32'hf309f4b7;
8'h51 : rvCrc[22] <= 32'hf545dd67;
8'h52 : rvCrc[22] <= 32'hff91a717;
8'h53 : rvCrc[22] <= 32'hf9dd8ec7;
8'h54 : rvCrc[22] <= 32'hea3953f7;
8'h55 : rvCrc[22] <= 32'hec757a27;
8'h56 : rvCrc[22] <= 32'he6a10057;
8'h57 : rvCrc[22] <= 32'he0ed2987;
8'h58 : rvCrc[22] <= 32'hc168ba37;
8'h59 : rvCrc[22] <= 32'hc72493e7;
8'h5a : rvCrc[22] <= 32'hcdf0e997;
8'h5b : rvCrc[22] <= 32'hcbbcc047;
8'h5c : rvCrc[22] <= 32'hd8581d77;
8'h5d : rvCrc[22] <= 32'hde1434a7;
8'h5e : rvCrc[22] <= 32'hd4c04ed7;
8'h5f : rvCrc[22] <= 32'hd28c6707;
8'h60 : rvCrc[22] <= 32'h5e4e53b7;
8'h61 : rvCrc[22] <= 32'h58027a67;
8'h62 : rvCrc[22] <= 32'h52d60017;
8'h63 : rvCrc[22] <= 32'h549a29c7;
8'h64 : rvCrc[22] <= 32'h477ef4f7;
8'h65 : rvCrc[22] <= 32'h4132dd27;
8'h66 : rvCrc[22] <= 32'h4be6a757;
8'h67 : rvCrc[22] <= 32'h4daa8e87;
8'h68 : rvCrc[22] <= 32'h6c2f1d37;
8'h69 : rvCrc[22] <= 32'h6a6334e7;
8'h6a : rvCrc[22] <= 32'h60b74e97;
8'h6b : rvCrc[22] <= 32'h66fb6747;
8'h6c : rvCrc[22] <= 32'h751fba77;
8'h6d : rvCrc[22] <= 32'h735393a7;
8'h6e : rvCrc[22] <= 32'h7987e9d7;
8'h6f : rvCrc[22] <= 32'h7fcbc007;
8'h70 : rvCrc[22] <= 32'h3a8cceb7;
8'h71 : rvCrc[22] <= 32'h3cc0e767;
8'h72 : rvCrc[22] <= 32'h36149d17;
8'h73 : rvCrc[22] <= 32'h3058b4c7;
8'h74 : rvCrc[22] <= 32'h23bc69f7;
8'h75 : rvCrc[22] <= 32'h25f04027;
8'h76 : rvCrc[22] <= 32'h2f243a57;
8'h77 : rvCrc[22] <= 32'h29681387;
8'h78 : rvCrc[22] <= 32'h08ed8037;
8'h79 : rvCrc[22] <= 32'h0ea1a9e7;
8'h7a : rvCrc[22] <= 32'h0475d397;
8'h7b : rvCrc[22] <= 32'h0239fa47;
8'h7c : rvCrc[22] <= 32'h11dd2777;
8'h7d : rvCrc[22] <= 32'h17910ea7;
8'h7e : rvCrc[22] <= 32'h1d4574d7;
8'h7f : rvCrc[22] <= 32'h1b095d07;
8'h80 : rvCrc[22] <= 32'h2b57ced9;
8'h81 : rvCrc[22] <= 32'h2d1be709;
8'h82 : rvCrc[22] <= 32'h27cf9d79;
8'h83 : rvCrc[22] <= 32'h2183b4a9;
8'h84 : rvCrc[22] <= 32'h32676999;
8'h85 : rvCrc[22] <= 32'h342b4049;
8'h86 : rvCrc[22] <= 32'h3eff3a39;
8'h87 : rvCrc[22] <= 32'h38b313e9;
8'h88 : rvCrc[22] <= 32'h19368059;
8'h89 : rvCrc[22] <= 32'h1f7aa989;
8'h8a : rvCrc[22] <= 32'h15aed3f9;
8'h8b : rvCrc[22] <= 32'h13e2fa29;
8'h8c : rvCrc[22] <= 32'h00062719;
8'h8d : rvCrc[22] <= 32'h064a0ec9;
8'h8e : rvCrc[22] <= 32'h0c9e74b9;
8'h8f : rvCrc[22] <= 32'h0ad25d69;
8'h90 : rvCrc[22] <= 32'h4f9553d9;
8'h91 : rvCrc[22] <= 32'h49d97a09;
8'h92 : rvCrc[22] <= 32'h430d0079;
8'h93 : rvCrc[22] <= 32'h454129a9;
8'h94 : rvCrc[22] <= 32'h56a5f499;
8'h95 : rvCrc[22] <= 32'h50e9dd49;
8'h96 : rvCrc[22] <= 32'h5a3da739;
8'h97 : rvCrc[22] <= 32'h5c718ee9;
8'h98 : rvCrc[22] <= 32'h7df41d59;
8'h99 : rvCrc[22] <= 32'h7bb83489;
8'h9a : rvCrc[22] <= 32'h716c4ef9;
8'h9b : rvCrc[22] <= 32'h77206729;
8'h9c : rvCrc[22] <= 32'h64c4ba19;
8'h9d : rvCrc[22] <= 32'h628893c9;
8'h9e : rvCrc[22] <= 32'h685ce9b9;
8'h9f : rvCrc[22] <= 32'h6e10c069;
8'ha0 : rvCrc[22] <= 32'he2d2f4d9;
8'ha1 : rvCrc[22] <= 32'he49edd09;
8'ha2 : rvCrc[22] <= 32'hee4aa779;
8'ha3 : rvCrc[22] <= 32'he8068ea9;
8'ha4 : rvCrc[22] <= 32'hfbe25399;
8'ha5 : rvCrc[22] <= 32'hfdae7a49;
8'ha6 : rvCrc[22] <= 32'hf77a0039;
8'ha7 : rvCrc[22] <= 32'hf13629e9;
8'ha8 : rvCrc[22] <= 32'hd0b3ba59;
8'ha9 : rvCrc[22] <= 32'hd6ff9389;
8'haa : rvCrc[22] <= 32'hdc2be9f9;
8'hab : rvCrc[22] <= 32'hda67c029;
8'hac : rvCrc[22] <= 32'hc9831d19;
8'had : rvCrc[22] <= 32'hcfcf34c9;
8'hae : rvCrc[22] <= 32'hc51b4eb9;
8'haf : rvCrc[22] <= 32'hc3576769;
8'hb0 : rvCrc[22] <= 32'h861069d9;
8'hb1 : rvCrc[22] <= 32'h805c4009;
8'hb2 : rvCrc[22] <= 32'h8a883a79;
8'hb3 : rvCrc[22] <= 32'h8cc413a9;
8'hb4 : rvCrc[22] <= 32'h9f20ce99;
8'hb5 : rvCrc[22] <= 32'h996ce749;
8'hb6 : rvCrc[22] <= 32'h93b89d39;
8'hb7 : rvCrc[22] <= 32'h95f4b4e9;
8'hb8 : rvCrc[22] <= 32'hb4712759;
8'hb9 : rvCrc[22] <= 32'hb23d0e89;
8'hba : rvCrc[22] <= 32'hb8e974f9;
8'hbb : rvCrc[22] <= 32'hbea55d29;
8'hbc : rvCrc[22] <= 32'had418019;
8'hbd : rvCrc[22] <= 32'hab0da9c9;
8'hbe : rvCrc[22] <= 32'ha1d9d3b9;
8'hbf : rvCrc[22] <= 32'ha795fa69;
8'hc0 : rvCrc[22] <= 32'hbc9ca76e;
8'hc1 : rvCrc[22] <= 32'hbad08ebe;
8'hc2 : rvCrc[22] <= 32'hb004f4ce;
8'hc3 : rvCrc[22] <= 32'hb648dd1e;
8'hc4 : rvCrc[22] <= 32'ha5ac002e;
8'hc5 : rvCrc[22] <= 32'ha3e029fe;
8'hc6 : rvCrc[22] <= 32'ha934538e;
8'hc7 : rvCrc[22] <= 32'haf787a5e;
8'hc8 : rvCrc[22] <= 32'h8efde9ee;
8'hc9 : rvCrc[22] <= 32'h88b1c03e;
8'hca : rvCrc[22] <= 32'h8265ba4e;
8'hcb : rvCrc[22] <= 32'h8429939e;
8'hcc : rvCrc[22] <= 32'h97cd4eae;
8'hcd : rvCrc[22] <= 32'h9181677e;
8'hce : rvCrc[22] <= 32'h9b551d0e;
8'hcf : rvCrc[22] <= 32'h9d1934de;
8'hd0 : rvCrc[22] <= 32'hd85e3a6e;
8'hd1 : rvCrc[22] <= 32'hde1213be;
8'hd2 : rvCrc[22] <= 32'hd4c669ce;
8'hd3 : rvCrc[22] <= 32'hd28a401e;
8'hd4 : rvCrc[22] <= 32'hc16e9d2e;
8'hd5 : rvCrc[22] <= 32'hc722b4fe;
8'hd6 : rvCrc[22] <= 32'hcdf6ce8e;
8'hd7 : rvCrc[22] <= 32'hcbbae75e;
8'hd8 : rvCrc[22] <= 32'hea3f74ee;
8'hd9 : rvCrc[22] <= 32'hec735d3e;
8'hda : rvCrc[22] <= 32'he6a7274e;
8'hdb : rvCrc[22] <= 32'he0eb0e9e;
8'hdc : rvCrc[22] <= 32'hf30fd3ae;
8'hdd : rvCrc[22] <= 32'hf543fa7e;
8'hde : rvCrc[22] <= 32'hff97800e;
8'hdf : rvCrc[22] <= 32'hf9dba9de;
8'he0 : rvCrc[22] <= 32'h75199d6e;
8'he1 : rvCrc[22] <= 32'h7355b4be;
8'he2 : rvCrc[22] <= 32'h7981cece;
8'he3 : rvCrc[22] <= 32'h7fcde71e;
8'he4 : rvCrc[22] <= 32'h6c293a2e;
8'he5 : rvCrc[22] <= 32'h6a6513fe;
8'he6 : rvCrc[22] <= 32'h60b1698e;
8'he7 : rvCrc[22] <= 32'h66fd405e;
8'he8 : rvCrc[22] <= 32'h4778d3ee;
8'he9 : rvCrc[22] <= 32'h4134fa3e;
8'hea : rvCrc[22] <= 32'h4be0804e;
8'heb : rvCrc[22] <= 32'h4daca99e;
8'hec : rvCrc[22] <= 32'h5e4874ae;
8'hed : rvCrc[22] <= 32'h58045d7e;
8'hee : rvCrc[22] <= 32'h52d0270e;
8'hef : rvCrc[22] <= 32'h549c0ede;
8'hf0 : rvCrc[22] <= 32'h11db006e;
8'hf1 : rvCrc[22] <= 32'h179729be;
8'hf2 : rvCrc[22] <= 32'h1d4353ce;
8'hf3 : rvCrc[22] <= 32'h1b0f7a1e;
8'hf4 : rvCrc[22] <= 32'h08eba72e;
8'hf5 : rvCrc[22] <= 32'h0ea78efe;
8'hf6 : rvCrc[22] <= 32'h0473f48e;
8'hf7 : rvCrc[22] <= 32'h023fdd5e;
8'hf8 : rvCrc[22] <= 32'h23ba4eee;
8'hf9 : rvCrc[22] <= 32'h25f6673e;
8'hfa : rvCrc[22] <= 32'h2f221d4e;
8'hfb : rvCrc[22] <= 32'h296e349e;
8'hfc : rvCrc[22] <= 32'h3a8ae9ae;
8'hfd : rvCrc[22] <= 32'h3cc6c07e;
8'hfe : rvCrc[22] <= 32'h3612ba0e;
8'hff : rvCrc[22] <= 32'h305e93de;
endcase
case(iv_Input[191:184])
8'h00 : rvCrc[23] <= 32'h00000000;
8'h01 : rvCrc[23] <= 32'h56af9db2;
8'h02 : rvCrc[23] <= 32'had5f3b64;
8'h03 : rvCrc[23] <= 32'hfbf0a6d6;
8'h04 : rvCrc[23] <= 32'h5e7f6b7f;
8'h05 : rvCrc[23] <= 32'h08d0f6cd;
8'h06 : rvCrc[23] <= 32'hf320501b;
8'h07 : rvCrc[23] <= 32'ha58fcda9;
8'h08 : rvCrc[23] <= 32'hbcfed6fe;
8'h09 : rvCrc[23] <= 32'hea514b4c;
8'h0a : rvCrc[23] <= 32'h11a1ed9a;
8'h0b : rvCrc[23] <= 32'h470e7028;
8'h0c : rvCrc[23] <= 32'he281bd81;
8'h0d : rvCrc[23] <= 32'hb42e2033;
8'h0e : rvCrc[23] <= 32'h4fde86e5;
8'h0f : rvCrc[23] <= 32'h19711b57;
8'h10 : rvCrc[23] <= 32'h7d3cb04b;
8'h11 : rvCrc[23] <= 32'h2b932df9;
8'h12 : rvCrc[23] <= 32'hd0638b2f;
8'h13 : rvCrc[23] <= 32'h86cc169d;
8'h14 : rvCrc[23] <= 32'h2343db34;
8'h15 : rvCrc[23] <= 32'h75ec4686;
8'h16 : rvCrc[23] <= 32'h8e1ce050;
8'h17 : rvCrc[23] <= 32'hd8b37de2;
8'h18 : rvCrc[23] <= 32'hc1c266b5;
8'h19 : rvCrc[23] <= 32'h976dfb07;
8'h1a : rvCrc[23] <= 32'h6c9d5dd1;
8'h1b : rvCrc[23] <= 32'h3a32c063;
8'h1c : rvCrc[23] <= 32'h9fbd0dca;
8'h1d : rvCrc[23] <= 32'hc9129078;
8'h1e : rvCrc[23] <= 32'h32e236ae;
8'h1f : rvCrc[23] <= 32'h644dab1c;
8'h20 : rvCrc[23] <= 32'hfa796096;
8'h21 : rvCrc[23] <= 32'hacd6fd24;
8'h22 : rvCrc[23] <= 32'h57265bf2;
8'h23 : rvCrc[23] <= 32'h0189c640;
8'h24 : rvCrc[23] <= 32'ha4060be9;
8'h25 : rvCrc[23] <= 32'hf2a9965b;
8'h26 : rvCrc[23] <= 32'h0959308d;
8'h27 : rvCrc[23] <= 32'h5ff6ad3f;
8'h28 : rvCrc[23] <= 32'h4687b668;
8'h29 : rvCrc[23] <= 32'h10282bda;
8'h2a : rvCrc[23] <= 32'hebd88d0c;
8'h2b : rvCrc[23] <= 32'hbd7710be;
8'h2c : rvCrc[23] <= 32'h18f8dd17;
8'h2d : rvCrc[23] <= 32'h4e5740a5;
8'h2e : rvCrc[23] <= 32'hb5a7e673;
8'h2f : rvCrc[23] <= 32'he3087bc1;
8'h30 : rvCrc[23] <= 32'h8745d0dd;
8'h31 : rvCrc[23] <= 32'hd1ea4d6f;
8'h32 : rvCrc[23] <= 32'h2a1aebb9;
8'h33 : rvCrc[23] <= 32'h7cb5760b;
8'h34 : rvCrc[23] <= 32'hd93abba2;
8'h35 : rvCrc[23] <= 32'h8f952610;
8'h36 : rvCrc[23] <= 32'h746580c6;
8'h37 : rvCrc[23] <= 32'h22ca1d74;
8'h38 : rvCrc[23] <= 32'h3bbb0623;
8'h39 : rvCrc[23] <= 32'h6d149b91;
8'h3a : rvCrc[23] <= 32'h96e43d47;
8'h3b : rvCrc[23] <= 32'hc04ba0f5;
8'h3c : rvCrc[23] <= 32'h65c46d5c;
8'h3d : rvCrc[23] <= 32'h336bf0ee;
8'h3e : rvCrc[23] <= 32'hc89b5638;
8'h3f : rvCrc[23] <= 32'h9e34cb8a;
8'h40 : rvCrc[23] <= 32'hf033dc9b;
8'h41 : rvCrc[23] <= 32'ha69c4129;
8'h42 : rvCrc[23] <= 32'h5d6ce7ff;
8'h43 : rvCrc[23] <= 32'h0bc37a4d;
8'h44 : rvCrc[23] <= 32'hae4cb7e4;
8'h45 : rvCrc[23] <= 32'hf8e32a56;
8'h46 : rvCrc[23] <= 32'h03138c80;
8'h47 : rvCrc[23] <= 32'h55bc1132;
8'h48 : rvCrc[23] <= 32'h4ccd0a65;
8'h49 : rvCrc[23] <= 32'h1a6297d7;
8'h4a : rvCrc[23] <= 32'he1923101;
8'h4b : rvCrc[23] <= 32'hb73dacb3;
8'h4c : rvCrc[23] <= 32'h12b2611a;
8'h4d : rvCrc[23] <= 32'h441dfca8;
8'h4e : rvCrc[23] <= 32'hbfed5a7e;
8'h4f : rvCrc[23] <= 32'he942c7cc;
8'h50 : rvCrc[23] <= 32'h8d0f6cd0;
8'h51 : rvCrc[23] <= 32'hdba0f162;
8'h52 : rvCrc[23] <= 32'h205057b4;
8'h53 : rvCrc[23] <= 32'h76ffca06;
8'h54 : rvCrc[23] <= 32'hd37007af;
8'h55 : rvCrc[23] <= 32'h85df9a1d;
8'h56 : rvCrc[23] <= 32'h7e2f3ccb;
8'h57 : rvCrc[23] <= 32'h2880a179;
8'h58 : rvCrc[23] <= 32'h31f1ba2e;
8'h59 : rvCrc[23] <= 32'h675e279c;
8'h5a : rvCrc[23] <= 32'h9cae814a;
8'h5b : rvCrc[23] <= 32'hca011cf8;
8'h5c : rvCrc[23] <= 32'h6f8ed151;
8'h5d : rvCrc[23] <= 32'h39214ce3;
8'h5e : rvCrc[23] <= 32'hc2d1ea35;
8'h5f : rvCrc[23] <= 32'h947e7787;
8'h60 : rvCrc[23] <= 32'h0a4abc0d;
8'h61 : rvCrc[23] <= 32'h5ce521bf;
8'h62 : rvCrc[23] <= 32'ha7158769;
8'h63 : rvCrc[23] <= 32'hf1ba1adb;
8'h64 : rvCrc[23] <= 32'h5435d772;
8'h65 : rvCrc[23] <= 32'h029a4ac0;
8'h66 : rvCrc[23] <= 32'hf96aec16;
8'h67 : rvCrc[23] <= 32'hafc571a4;
8'h68 : rvCrc[23] <= 32'hb6b46af3;
8'h69 : rvCrc[23] <= 32'he01bf741;
8'h6a : rvCrc[23] <= 32'h1beb5197;
8'h6b : rvCrc[23] <= 32'h4d44cc25;
8'h6c : rvCrc[23] <= 32'he8cb018c;
8'h6d : rvCrc[23] <= 32'hbe649c3e;
8'h6e : rvCrc[23] <= 32'h45943ae8;
8'h6f : rvCrc[23] <= 32'h133ba75a;
8'h70 : rvCrc[23] <= 32'h77760c46;
8'h71 : rvCrc[23] <= 32'h21d991f4;
8'h72 : rvCrc[23] <= 32'hda293722;
8'h73 : rvCrc[23] <= 32'h8c86aa90;
8'h74 : rvCrc[23] <= 32'h29096739;
8'h75 : rvCrc[23] <= 32'h7fa6fa8b;
8'h76 : rvCrc[23] <= 32'h84565c5d;
8'h77 : rvCrc[23] <= 32'hd2f9c1ef;
8'h78 : rvCrc[23] <= 32'hcb88dab8;
8'h79 : rvCrc[23] <= 32'h9d27470a;
8'h7a : rvCrc[23] <= 32'h66d7e1dc;
8'h7b : rvCrc[23] <= 32'h30787c6e;
8'h7c : rvCrc[23] <= 32'h95f7b1c7;
8'h7d : rvCrc[23] <= 32'hc3582c75;
8'h7e : rvCrc[23] <= 32'h38a88aa3;
8'h7f : rvCrc[23] <= 32'h6e071711;
8'h80 : rvCrc[23] <= 32'he4a6a481;
8'h81 : rvCrc[23] <= 32'hb2093933;
8'h82 : rvCrc[23] <= 32'h49f99fe5;
8'h83 : rvCrc[23] <= 32'h1f560257;
8'h84 : rvCrc[23] <= 32'hbad9cffe;
8'h85 : rvCrc[23] <= 32'hec76524c;
8'h86 : rvCrc[23] <= 32'h1786f49a;
8'h87 : rvCrc[23] <= 32'h41296928;
8'h88 : rvCrc[23] <= 32'h5858727f;
8'h89 : rvCrc[23] <= 32'h0ef7efcd;
8'h8a : rvCrc[23] <= 32'hf507491b;
8'h8b : rvCrc[23] <= 32'ha3a8d4a9;
8'h8c : rvCrc[23] <= 32'h06271900;
8'h8d : rvCrc[23] <= 32'h508884b2;
8'h8e : rvCrc[23] <= 32'hab782264;
8'h8f : rvCrc[23] <= 32'hfdd7bfd6;
8'h90 : rvCrc[23] <= 32'h999a14ca;
8'h91 : rvCrc[23] <= 32'hcf358978;
8'h92 : rvCrc[23] <= 32'h34c52fae;
8'h93 : rvCrc[23] <= 32'h626ab21c;
8'h94 : rvCrc[23] <= 32'hc7e57fb5;
8'h95 : rvCrc[23] <= 32'h914ae207;
8'h96 : rvCrc[23] <= 32'h6aba44d1;
8'h97 : rvCrc[23] <= 32'h3c15d963;
8'h98 : rvCrc[23] <= 32'h2564c234;
8'h99 : rvCrc[23] <= 32'h73cb5f86;
8'h9a : rvCrc[23] <= 32'h883bf950;
8'h9b : rvCrc[23] <= 32'hde9464e2;
8'h9c : rvCrc[23] <= 32'h7b1ba94b;
8'h9d : rvCrc[23] <= 32'h2db434f9;
8'h9e : rvCrc[23] <= 32'hd644922f;
8'h9f : rvCrc[23] <= 32'h80eb0f9d;
8'ha0 : rvCrc[23] <= 32'h1edfc417;
8'ha1 : rvCrc[23] <= 32'h487059a5;
8'ha2 : rvCrc[23] <= 32'hb380ff73;
8'ha3 : rvCrc[23] <= 32'he52f62c1;
8'ha4 : rvCrc[23] <= 32'h40a0af68;
8'ha5 : rvCrc[23] <= 32'h160f32da;
8'ha6 : rvCrc[23] <= 32'hedff940c;
8'ha7 : rvCrc[23] <= 32'hbb5009be;
8'ha8 : rvCrc[23] <= 32'ha22112e9;
8'ha9 : rvCrc[23] <= 32'hf48e8f5b;
8'haa : rvCrc[23] <= 32'h0f7e298d;
8'hab : rvCrc[23] <= 32'h59d1b43f;
8'hac : rvCrc[23] <= 32'hfc5e7996;
8'had : rvCrc[23] <= 32'haaf1e424;
8'hae : rvCrc[23] <= 32'h510142f2;
8'haf : rvCrc[23] <= 32'h07aedf40;
8'hb0 : rvCrc[23] <= 32'h63e3745c;
8'hb1 : rvCrc[23] <= 32'h354ce9ee;
8'hb2 : rvCrc[23] <= 32'hcebc4f38;
8'hb3 : rvCrc[23] <= 32'h9813d28a;
8'hb4 : rvCrc[23] <= 32'h3d9c1f23;
8'hb5 : rvCrc[23] <= 32'h6b338291;
8'hb6 : rvCrc[23] <= 32'h90c32447;
8'hb7 : rvCrc[23] <= 32'hc66cb9f5;
8'hb8 : rvCrc[23] <= 32'hdf1da2a2;
8'hb9 : rvCrc[23] <= 32'h89b23f10;
8'hba : rvCrc[23] <= 32'h724299c6;
8'hbb : rvCrc[23] <= 32'h24ed0474;
8'hbc : rvCrc[23] <= 32'h8162c9dd;
8'hbd : rvCrc[23] <= 32'hd7cd546f;
8'hbe : rvCrc[23] <= 32'h2c3df2b9;
8'hbf : rvCrc[23] <= 32'h7a926f0b;
8'hc0 : rvCrc[23] <= 32'h1495781a;
8'hc1 : rvCrc[23] <= 32'h423ae5a8;
8'hc2 : rvCrc[23] <= 32'hb9ca437e;
8'hc3 : rvCrc[23] <= 32'hef65decc;
8'hc4 : rvCrc[23] <= 32'h4aea1365;
8'hc5 : rvCrc[23] <= 32'h1c458ed7;
8'hc6 : rvCrc[23] <= 32'he7b52801;
8'hc7 : rvCrc[23] <= 32'hb11ab5b3;
8'hc8 : rvCrc[23] <= 32'ha86baee4;
8'hc9 : rvCrc[23] <= 32'hfec43356;
8'hca : rvCrc[23] <= 32'h05349580;
8'hcb : rvCrc[23] <= 32'h539b0832;
8'hcc : rvCrc[23] <= 32'hf614c59b;
8'hcd : rvCrc[23] <= 32'ha0bb5829;
8'hce : rvCrc[23] <= 32'h5b4bfeff;
8'hcf : rvCrc[23] <= 32'h0de4634d;
8'hd0 : rvCrc[23] <= 32'h69a9c851;
8'hd1 : rvCrc[23] <= 32'h3f0655e3;
8'hd2 : rvCrc[23] <= 32'hc4f6f335;
8'hd3 : rvCrc[23] <= 32'h92596e87;
8'hd4 : rvCrc[23] <= 32'h37d6a32e;
8'hd5 : rvCrc[23] <= 32'h61793e9c;
8'hd6 : rvCrc[23] <= 32'h9a89984a;
8'hd7 : rvCrc[23] <= 32'hcc2605f8;
8'hd8 : rvCrc[23] <= 32'hd5571eaf;
8'hd9 : rvCrc[23] <= 32'h83f8831d;
8'hda : rvCrc[23] <= 32'h780825cb;
8'hdb : rvCrc[23] <= 32'h2ea7b879;
8'hdc : rvCrc[23] <= 32'h8b2875d0;
8'hdd : rvCrc[23] <= 32'hdd87e862;
8'hde : rvCrc[23] <= 32'h26774eb4;
8'hdf : rvCrc[23] <= 32'h70d8d306;
8'he0 : rvCrc[23] <= 32'heeec188c;
8'he1 : rvCrc[23] <= 32'hb843853e;
8'he2 : rvCrc[23] <= 32'h43b323e8;
8'he3 : rvCrc[23] <= 32'h151cbe5a;
8'he4 : rvCrc[23] <= 32'hb09373f3;
8'he5 : rvCrc[23] <= 32'he63cee41;
8'he6 : rvCrc[23] <= 32'h1dcc4897;
8'he7 : rvCrc[23] <= 32'h4b63d525;
8'he8 : rvCrc[23] <= 32'h5212ce72;
8'he9 : rvCrc[23] <= 32'h04bd53c0;
8'hea : rvCrc[23] <= 32'hff4df516;
8'heb : rvCrc[23] <= 32'ha9e268a4;
8'hec : rvCrc[23] <= 32'h0c6da50d;
8'hed : rvCrc[23] <= 32'h5ac238bf;
8'hee : rvCrc[23] <= 32'ha1329e69;
8'hef : rvCrc[23] <= 32'hf79d03db;
8'hf0 : rvCrc[23] <= 32'h93d0a8c7;
8'hf1 : rvCrc[23] <= 32'hc57f3575;
8'hf2 : rvCrc[23] <= 32'h3e8f93a3;
8'hf3 : rvCrc[23] <= 32'h68200e11;
8'hf4 : rvCrc[23] <= 32'hcdafc3b8;
8'hf5 : rvCrc[23] <= 32'h9b005e0a;
8'hf6 : rvCrc[23] <= 32'h60f0f8dc;
8'hf7 : rvCrc[23] <= 32'h365f656e;
8'hf8 : rvCrc[23] <= 32'h2f2e7e39;
8'hf9 : rvCrc[23] <= 32'h7981e38b;
8'hfa : rvCrc[23] <= 32'h8271455d;
8'hfb : rvCrc[23] <= 32'hd4ded8ef;
8'hfc : rvCrc[23] <= 32'h71511546;
8'hfd : rvCrc[23] <= 32'h27fe88f4;
8'hfe : rvCrc[23] <= 32'hdc0e2e22;
8'hff : rvCrc[23] <= 32'h8aa1b390;
endcase
case(iv_Input[199:192])
8'h00 : rvCrc[24] <= 32'h00000000;
8'h01 : rvCrc[24] <= 32'hcd8c54b5;
8'h02 : rvCrc[24] <= 32'h9fd9b4dd;
8'h03 : rvCrc[24] <= 32'h5255e068;
8'h04 : rvCrc[24] <= 32'h3b72740d;
8'h05 : rvCrc[24] <= 32'hf6fe20b8;
8'h06 : rvCrc[24] <= 32'ha4abc0d0;
8'h07 : rvCrc[24] <= 32'h69279465;
8'h08 : rvCrc[24] <= 32'h76e4e81a;
8'h09 : rvCrc[24] <= 32'hbb68bcaf;
8'h0a : rvCrc[24] <= 32'he93d5cc7;
8'h0b : rvCrc[24] <= 32'h24b10872;
8'h0c : rvCrc[24] <= 32'h4d969c17;
8'h0d : rvCrc[24] <= 32'h801ac8a2;
8'h0e : rvCrc[24] <= 32'hd24f28ca;
8'h0f : rvCrc[24] <= 32'h1fc37c7f;
8'h10 : rvCrc[24] <= 32'hedc9d034;
8'h11 : rvCrc[24] <= 32'h20458481;
8'h12 : rvCrc[24] <= 32'h721064e9;
8'h13 : rvCrc[24] <= 32'hbf9c305c;
8'h14 : rvCrc[24] <= 32'hd6bba439;
8'h15 : rvCrc[24] <= 32'h1b37f08c;
8'h16 : rvCrc[24] <= 32'h496210e4;
8'h17 : rvCrc[24] <= 32'h84ee4451;
8'h18 : rvCrc[24] <= 32'h9b2d382e;
8'h19 : rvCrc[24] <= 32'h56a16c9b;
8'h1a : rvCrc[24] <= 32'h04f48cf3;
8'h1b : rvCrc[24] <= 32'hc978d846;
8'h1c : rvCrc[24] <= 32'ha05f4c23;
8'h1d : rvCrc[24] <= 32'h6dd31896;
8'h1e : rvCrc[24] <= 32'h3f86f8fe;
8'h1f : rvCrc[24] <= 32'hf20aac4b;
8'h20 : rvCrc[24] <= 32'hdf52bddf;
8'h21 : rvCrc[24] <= 32'h12dee96a;
8'h22 : rvCrc[24] <= 32'h408b0902;
8'h23 : rvCrc[24] <= 32'h8d075db7;
8'h24 : rvCrc[24] <= 32'he420c9d2;
8'h25 : rvCrc[24] <= 32'h29ac9d67;
8'h26 : rvCrc[24] <= 32'h7bf97d0f;
8'h27 : rvCrc[24] <= 32'hb67529ba;
8'h28 : rvCrc[24] <= 32'ha9b655c5;
8'h29 : rvCrc[24] <= 32'h643a0170;
8'h2a : rvCrc[24] <= 32'h366fe118;
8'h2b : rvCrc[24] <= 32'hfbe3b5ad;
8'h2c : rvCrc[24] <= 32'h92c421c8;
8'h2d : rvCrc[24] <= 32'h5f48757d;
8'h2e : rvCrc[24] <= 32'h0d1d9515;
8'h2f : rvCrc[24] <= 32'hc091c1a0;
8'h30 : rvCrc[24] <= 32'h329b6deb;
8'h31 : rvCrc[24] <= 32'hff17395e;
8'h32 : rvCrc[24] <= 32'had42d936;
8'h33 : rvCrc[24] <= 32'h60ce8d83;
8'h34 : rvCrc[24] <= 32'h09e919e6;
8'h35 : rvCrc[24] <= 32'hc4654d53;
8'h36 : rvCrc[24] <= 32'h9630ad3b;
8'h37 : rvCrc[24] <= 32'h5bbcf98e;
8'h38 : rvCrc[24] <= 32'h447f85f1;
8'h39 : rvCrc[24] <= 32'h89f3d144;
8'h3a : rvCrc[24] <= 32'hdba6312c;
8'h3b : rvCrc[24] <= 32'h162a6599;
8'h3c : rvCrc[24] <= 32'h7f0df1fc;
8'h3d : rvCrc[24] <= 32'hb281a549;
8'h3e : rvCrc[24] <= 32'he0d44521;
8'h3f : rvCrc[24] <= 32'h2d581194;
8'h40 : rvCrc[24] <= 32'hba646609;
8'h41 : rvCrc[24] <= 32'h77e832bc;
8'h42 : rvCrc[24] <= 32'h25bdd2d4;
8'h43 : rvCrc[24] <= 32'he8318661;
8'h44 : rvCrc[24] <= 32'h81161204;
8'h45 : rvCrc[24] <= 32'h4c9a46b1;
8'h46 : rvCrc[24] <= 32'h1ecfa6d9;
8'h47 : rvCrc[24] <= 32'hd343f26c;
8'h48 : rvCrc[24] <= 32'hcc808e13;
8'h49 : rvCrc[24] <= 32'h010cdaa6;
8'h4a : rvCrc[24] <= 32'h53593ace;
8'h4b : rvCrc[24] <= 32'h9ed56e7b;
8'h4c : rvCrc[24] <= 32'hf7f2fa1e;
8'h4d : rvCrc[24] <= 32'h3a7eaeab;
8'h4e : rvCrc[24] <= 32'h682b4ec3;
8'h4f : rvCrc[24] <= 32'ha5a71a76;
8'h50 : rvCrc[24] <= 32'h57adb63d;
8'h51 : rvCrc[24] <= 32'h9a21e288;
8'h52 : rvCrc[24] <= 32'hc87402e0;
8'h53 : rvCrc[24] <= 32'h05f85655;
8'h54 : rvCrc[24] <= 32'h6cdfc230;
8'h55 : rvCrc[24] <= 32'ha1539685;
8'h56 : rvCrc[24] <= 32'hf30676ed;
8'h57 : rvCrc[24] <= 32'h3e8a2258;
8'h58 : rvCrc[24] <= 32'h21495e27;
8'h59 : rvCrc[24] <= 32'hecc50a92;
8'h5a : rvCrc[24] <= 32'hbe90eafa;
8'h5b : rvCrc[24] <= 32'h731cbe4f;
8'h5c : rvCrc[24] <= 32'h1a3b2a2a;
8'h5d : rvCrc[24] <= 32'hd7b77e9f;
8'h5e : rvCrc[24] <= 32'h85e29ef7;
8'h5f : rvCrc[24] <= 32'h486eca42;
8'h60 : rvCrc[24] <= 32'h6536dbd6;
8'h61 : rvCrc[24] <= 32'ha8ba8f63;
8'h62 : rvCrc[24] <= 32'hfaef6f0b;
8'h63 : rvCrc[24] <= 32'h37633bbe;
8'h64 : rvCrc[24] <= 32'h5e44afdb;
8'h65 : rvCrc[24] <= 32'h93c8fb6e;
8'h66 : rvCrc[24] <= 32'hc19d1b06;
8'h67 : rvCrc[24] <= 32'h0c114fb3;
8'h68 : rvCrc[24] <= 32'h13d233cc;
8'h69 : rvCrc[24] <= 32'hde5e6779;
8'h6a : rvCrc[24] <= 32'h8c0b8711;
8'h6b : rvCrc[24] <= 32'h4187d3a4;
8'h6c : rvCrc[24] <= 32'h28a047c1;
8'h6d : rvCrc[24] <= 32'he52c1374;
8'h6e : rvCrc[24] <= 32'hb779f31c;
8'h6f : rvCrc[24] <= 32'h7af5a7a9;
8'h70 : rvCrc[24] <= 32'h88ff0be2;
8'h71 : rvCrc[24] <= 32'h45735f57;
8'h72 : rvCrc[24] <= 32'h1726bf3f;
8'h73 : rvCrc[24] <= 32'hdaaaeb8a;
8'h74 : rvCrc[24] <= 32'hb38d7fef;
8'h75 : rvCrc[24] <= 32'h7e012b5a;
8'h76 : rvCrc[24] <= 32'h2c54cb32;
8'h77 : rvCrc[24] <= 32'he1d89f87;
8'h78 : rvCrc[24] <= 32'hfe1be3f8;
8'h79 : rvCrc[24] <= 32'h3397b74d;
8'h7a : rvCrc[24] <= 32'h61c25725;
8'h7b : rvCrc[24] <= 32'hac4e0390;
8'h7c : rvCrc[24] <= 32'hc56997f5;
8'h7d : rvCrc[24] <= 32'h08e5c340;
8'h7e : rvCrc[24] <= 32'h5ab02328;
8'h7f : rvCrc[24] <= 32'h973c779d;
8'h80 : rvCrc[24] <= 32'h7009d1a5;
8'h81 : rvCrc[24] <= 32'hbd858510;
8'h82 : rvCrc[24] <= 32'hefd06578;
8'h83 : rvCrc[24] <= 32'h225c31cd;
8'h84 : rvCrc[24] <= 32'h4b7ba5a8;
8'h85 : rvCrc[24] <= 32'h86f7f11d;
8'h86 : rvCrc[24] <= 32'hd4a21175;
8'h87 : rvCrc[24] <= 32'h192e45c0;
8'h88 : rvCrc[24] <= 32'h06ed39bf;
8'h89 : rvCrc[24] <= 32'hcb616d0a;
8'h8a : rvCrc[24] <= 32'h99348d62;
8'h8b : rvCrc[24] <= 32'h54b8d9d7;
8'h8c : rvCrc[24] <= 32'h3d9f4db2;
8'h8d : rvCrc[24] <= 32'hf0131907;
8'h8e : rvCrc[24] <= 32'ha246f96f;
8'h8f : rvCrc[24] <= 32'h6fcaadda;
8'h90 : rvCrc[24] <= 32'h9dc00191;
8'h91 : rvCrc[24] <= 32'h504c5524;
8'h92 : rvCrc[24] <= 32'h0219b54c;
8'h93 : rvCrc[24] <= 32'hcf95e1f9;
8'h94 : rvCrc[24] <= 32'ha6b2759c;
8'h95 : rvCrc[24] <= 32'h6b3e2129;
8'h96 : rvCrc[24] <= 32'h396bc141;
8'h97 : rvCrc[24] <= 32'hf4e795f4;
8'h98 : rvCrc[24] <= 32'heb24e98b;
8'h99 : rvCrc[24] <= 32'h26a8bd3e;
8'h9a : rvCrc[24] <= 32'h74fd5d56;
8'h9b : rvCrc[24] <= 32'hb97109e3;
8'h9c : rvCrc[24] <= 32'hd0569d86;
8'h9d : rvCrc[24] <= 32'h1ddac933;
8'h9e : rvCrc[24] <= 32'h4f8f295b;
8'h9f : rvCrc[24] <= 32'h82037dee;
8'ha0 : rvCrc[24] <= 32'haf5b6c7a;
8'ha1 : rvCrc[24] <= 32'h62d738cf;
8'ha2 : rvCrc[24] <= 32'h3082d8a7;
8'ha3 : rvCrc[24] <= 32'hfd0e8c12;
8'ha4 : rvCrc[24] <= 32'h94291877;
8'ha5 : rvCrc[24] <= 32'h59a54cc2;
8'ha6 : rvCrc[24] <= 32'h0bf0acaa;
8'ha7 : rvCrc[24] <= 32'hc67cf81f;
8'ha8 : rvCrc[24] <= 32'hd9bf8460;
8'ha9 : rvCrc[24] <= 32'h1433d0d5;
8'haa : rvCrc[24] <= 32'h466630bd;
8'hab : rvCrc[24] <= 32'h8bea6408;
8'hac : rvCrc[24] <= 32'he2cdf06d;
8'had : rvCrc[24] <= 32'h2f41a4d8;
8'hae : rvCrc[24] <= 32'h7d1444b0;
8'haf : rvCrc[24] <= 32'hb0981005;
8'hb0 : rvCrc[24] <= 32'h4292bc4e;
8'hb1 : rvCrc[24] <= 32'h8f1ee8fb;
8'hb2 : rvCrc[24] <= 32'hdd4b0893;
8'hb3 : rvCrc[24] <= 32'h10c75c26;
8'hb4 : rvCrc[24] <= 32'h79e0c843;
8'hb5 : rvCrc[24] <= 32'hb46c9cf6;
8'hb6 : rvCrc[24] <= 32'he6397c9e;
8'hb7 : rvCrc[24] <= 32'h2bb5282b;
8'hb8 : rvCrc[24] <= 32'h34765454;
8'hb9 : rvCrc[24] <= 32'hf9fa00e1;
8'hba : rvCrc[24] <= 32'habafe089;
8'hbb : rvCrc[24] <= 32'h6623b43c;
8'hbc : rvCrc[24] <= 32'h0f042059;
8'hbd : rvCrc[24] <= 32'hc28874ec;
8'hbe : rvCrc[24] <= 32'h90dd9484;
8'hbf : rvCrc[24] <= 32'h5d51c031;
8'hc0 : rvCrc[24] <= 32'hca6db7ac;
8'hc1 : rvCrc[24] <= 32'h07e1e319;
8'hc2 : rvCrc[24] <= 32'h55b40371;
8'hc3 : rvCrc[24] <= 32'h983857c4;
8'hc4 : rvCrc[24] <= 32'hf11fc3a1;
8'hc5 : rvCrc[24] <= 32'h3c939714;
8'hc6 : rvCrc[24] <= 32'h6ec6777c;
8'hc7 : rvCrc[24] <= 32'ha34a23c9;
8'hc8 : rvCrc[24] <= 32'hbc895fb6;
8'hc9 : rvCrc[24] <= 32'h71050b03;
8'hca : rvCrc[24] <= 32'h2350eb6b;
8'hcb : rvCrc[24] <= 32'heedcbfde;
8'hcc : rvCrc[24] <= 32'h87fb2bbb;
8'hcd : rvCrc[24] <= 32'h4a777f0e;
8'hce : rvCrc[24] <= 32'h18229f66;
8'hcf : rvCrc[24] <= 32'hd5aecbd3;
8'hd0 : rvCrc[24] <= 32'h27a46798;
8'hd1 : rvCrc[24] <= 32'hea28332d;
8'hd2 : rvCrc[24] <= 32'hb87dd345;
8'hd3 : rvCrc[24] <= 32'h75f187f0;
8'hd4 : rvCrc[24] <= 32'h1cd61395;
8'hd5 : rvCrc[24] <= 32'hd15a4720;
8'hd6 : rvCrc[24] <= 32'h830fa748;
8'hd7 : rvCrc[24] <= 32'h4e83f3fd;
8'hd8 : rvCrc[24] <= 32'h51408f82;
8'hd9 : rvCrc[24] <= 32'h9cccdb37;
8'hda : rvCrc[24] <= 32'hce993b5f;
8'hdb : rvCrc[24] <= 32'h03156fea;
8'hdc : rvCrc[24] <= 32'h6a32fb8f;
8'hdd : rvCrc[24] <= 32'ha7beaf3a;
8'hde : rvCrc[24] <= 32'hf5eb4f52;
8'hdf : rvCrc[24] <= 32'h38671be7;
8'he0 : rvCrc[24] <= 32'h153f0a73;
8'he1 : rvCrc[24] <= 32'hd8b35ec6;
8'he2 : rvCrc[24] <= 32'h8ae6beae;
8'he3 : rvCrc[24] <= 32'h476aea1b;
8'he4 : rvCrc[24] <= 32'h2e4d7e7e;
8'he5 : rvCrc[24] <= 32'he3c12acb;
8'he6 : rvCrc[24] <= 32'hb194caa3;
8'he7 : rvCrc[24] <= 32'h7c189e16;
8'he8 : rvCrc[24] <= 32'h63dbe269;
8'he9 : rvCrc[24] <= 32'hae57b6dc;
8'hea : rvCrc[24] <= 32'hfc0256b4;
8'heb : rvCrc[24] <= 32'h318e0201;
8'hec : rvCrc[24] <= 32'h58a99664;
8'hed : rvCrc[24] <= 32'h9525c2d1;
8'hee : rvCrc[24] <= 32'hc77022b9;
8'hef : rvCrc[24] <= 32'h0afc760c;
8'hf0 : rvCrc[24] <= 32'hf8f6da47;
8'hf1 : rvCrc[24] <= 32'h357a8ef2;
8'hf2 : rvCrc[24] <= 32'h672f6e9a;
8'hf3 : rvCrc[24] <= 32'haaa33a2f;
8'hf4 : rvCrc[24] <= 32'hc384ae4a;
8'hf5 : rvCrc[24] <= 32'h0e08faff;
8'hf6 : rvCrc[24] <= 32'h5c5d1a97;
8'hf7 : rvCrc[24] <= 32'h91d14e22;
8'hf8 : rvCrc[24] <= 32'h8e12325d;
8'hf9 : rvCrc[24] <= 32'h439e66e8;
8'hfa : rvCrc[24] <= 32'h11cb8680;
8'hfb : rvCrc[24] <= 32'hdc47d235;
8'hfc : rvCrc[24] <= 32'hb5604650;
8'hfd : rvCrc[24] <= 32'h78ec12e5;
8'hfe : rvCrc[24] <= 32'h2ab9f28d;
8'hff : rvCrc[24] <= 32'he735a638;
endcase
case(iv_Input[207:200])
8'h00 : rvCrc[25] <= 32'h00000000;
8'h01 : rvCrc[25] <= 32'he013a34a;
8'h02 : rvCrc[25] <= 32'hc4e65b23;
8'h03 : rvCrc[25] <= 32'h24f5f869;
8'h04 : rvCrc[25] <= 32'h8d0dabf1;
8'h05 : rvCrc[25] <= 32'h6d1e08bb;
8'h06 : rvCrc[25] <= 32'h49ebf0d2;
8'h07 : rvCrc[25] <= 32'ha9f85398;
8'h08 : rvCrc[25] <= 32'h1eda4a55;
8'h09 : rvCrc[25] <= 32'hfec9e91f;
8'h0a : rvCrc[25] <= 32'hda3c1176;
8'h0b : rvCrc[25] <= 32'h3a2fb23c;
8'h0c : rvCrc[25] <= 32'h93d7e1a4;
8'h0d : rvCrc[25] <= 32'h73c442ee;
8'h0e : rvCrc[25] <= 32'h5731ba87;
8'h0f : rvCrc[25] <= 32'hb72219cd;
8'h10 : rvCrc[25] <= 32'h3db494aa;
8'h11 : rvCrc[25] <= 32'hdda737e0;
8'h12 : rvCrc[25] <= 32'hf952cf89;
8'h13 : rvCrc[25] <= 32'h19416cc3;
8'h14 : rvCrc[25] <= 32'hb0b93f5b;
8'h15 : rvCrc[25] <= 32'h50aa9c11;
8'h16 : rvCrc[25] <= 32'h745f6478;
8'h17 : rvCrc[25] <= 32'h944cc732;
8'h18 : rvCrc[25] <= 32'h236edeff;
8'h19 : rvCrc[25] <= 32'hc37d7db5;
8'h1a : rvCrc[25] <= 32'he78885dc;
8'h1b : rvCrc[25] <= 32'h079b2696;
8'h1c : rvCrc[25] <= 32'hae63750e;
8'h1d : rvCrc[25] <= 32'h4e70d644;
8'h1e : rvCrc[25] <= 32'h6a852e2d;
8'h1f : rvCrc[25] <= 32'h8a968d67;
8'h20 : rvCrc[25] <= 32'h7b692954;
8'h21 : rvCrc[25] <= 32'h9b7a8a1e;
8'h22 : rvCrc[25] <= 32'hbf8f7277;
8'h23 : rvCrc[25] <= 32'h5f9cd13d;
8'h24 : rvCrc[25] <= 32'hf66482a5;
8'h25 : rvCrc[25] <= 32'h167721ef;
8'h26 : rvCrc[25] <= 32'h3282d986;
8'h27 : rvCrc[25] <= 32'hd2917acc;
8'h28 : rvCrc[25] <= 32'h65b36301;
8'h29 : rvCrc[25] <= 32'h85a0c04b;
8'h2a : rvCrc[25] <= 32'ha1553822;
8'h2b : rvCrc[25] <= 32'h41469b68;
8'h2c : rvCrc[25] <= 32'he8bec8f0;
8'h2d : rvCrc[25] <= 32'h08ad6bba;
8'h2e : rvCrc[25] <= 32'h2c5893d3;
8'h2f : rvCrc[25] <= 32'hcc4b3099;
8'h30 : rvCrc[25] <= 32'h46ddbdfe;
8'h31 : rvCrc[25] <= 32'ha6ce1eb4;
8'h32 : rvCrc[25] <= 32'h823be6dd;
8'h33 : rvCrc[25] <= 32'h62284597;
8'h34 : rvCrc[25] <= 32'hcbd0160f;
8'h35 : rvCrc[25] <= 32'h2bc3b545;
8'h36 : rvCrc[25] <= 32'h0f364d2c;
8'h37 : rvCrc[25] <= 32'hef25ee66;
8'h38 : rvCrc[25] <= 32'h5807f7ab;
8'h39 : rvCrc[25] <= 32'hb81454e1;
8'h3a : rvCrc[25] <= 32'h9ce1ac88;
8'h3b : rvCrc[25] <= 32'h7cf20fc2;
8'h3c : rvCrc[25] <= 32'hd50a5c5a;
8'h3d : rvCrc[25] <= 32'h3519ff10;
8'h3e : rvCrc[25] <= 32'h11ec0779;
8'h3f : rvCrc[25] <= 32'hf1ffa433;
8'h40 : rvCrc[25] <= 32'hf6d252a8;
8'h41 : rvCrc[25] <= 32'h16c1f1e2;
8'h42 : rvCrc[25] <= 32'h3234098b;
8'h43 : rvCrc[25] <= 32'hd227aac1;
8'h44 : rvCrc[25] <= 32'h7bdff959;
8'h45 : rvCrc[25] <= 32'h9bcc5a13;
8'h46 : rvCrc[25] <= 32'hbf39a27a;
8'h47 : rvCrc[25] <= 32'h5f2a0130;
8'h48 : rvCrc[25] <= 32'he80818fd;
8'h49 : rvCrc[25] <= 32'h081bbbb7;
8'h4a : rvCrc[25] <= 32'h2cee43de;
8'h4b : rvCrc[25] <= 32'hccfde094;
8'h4c : rvCrc[25] <= 32'h6505b30c;
8'h4d : rvCrc[25] <= 32'h85161046;
8'h4e : rvCrc[25] <= 32'ha1e3e82f;
8'h4f : rvCrc[25] <= 32'h41f04b65;
8'h50 : rvCrc[25] <= 32'hcb66c602;
8'h51 : rvCrc[25] <= 32'h2b756548;
8'h52 : rvCrc[25] <= 32'h0f809d21;
8'h53 : rvCrc[25] <= 32'hef933e6b;
8'h54 : rvCrc[25] <= 32'h466b6df3;
8'h55 : rvCrc[25] <= 32'ha678ceb9;
8'h56 : rvCrc[25] <= 32'h828d36d0;
8'h57 : rvCrc[25] <= 32'h629e959a;
8'h58 : rvCrc[25] <= 32'hd5bc8c57;
8'h59 : rvCrc[25] <= 32'h35af2f1d;
8'h5a : rvCrc[25] <= 32'h115ad774;
8'h5b : rvCrc[25] <= 32'hf149743e;
8'h5c : rvCrc[25] <= 32'h58b127a6;
8'h5d : rvCrc[25] <= 32'hb8a284ec;
8'h5e : rvCrc[25] <= 32'h9c577c85;
8'h5f : rvCrc[25] <= 32'h7c44dfcf;
8'h60 : rvCrc[25] <= 32'h8dbb7bfc;
8'h61 : rvCrc[25] <= 32'h6da8d8b6;
8'h62 : rvCrc[25] <= 32'h495d20df;
8'h63 : rvCrc[25] <= 32'ha94e8395;
8'h64 : rvCrc[25] <= 32'h00b6d00d;
8'h65 : rvCrc[25] <= 32'he0a57347;
8'h66 : rvCrc[25] <= 32'hc4508b2e;
8'h67 : rvCrc[25] <= 32'h24432864;
8'h68 : rvCrc[25] <= 32'h936131a9;
8'h69 : rvCrc[25] <= 32'h737292e3;
8'h6a : rvCrc[25] <= 32'h57876a8a;
8'h6b : rvCrc[25] <= 32'hb794c9c0;
8'h6c : rvCrc[25] <= 32'h1e6c9a58;
8'h6d : rvCrc[25] <= 32'hfe7f3912;
8'h6e : rvCrc[25] <= 32'hda8ac17b;
8'h6f : rvCrc[25] <= 32'h3a996231;
8'h70 : rvCrc[25] <= 32'hb00fef56;
8'h71 : rvCrc[25] <= 32'h501c4c1c;
8'h72 : rvCrc[25] <= 32'h74e9b475;
8'h73 : rvCrc[25] <= 32'h94fa173f;
8'h74 : rvCrc[25] <= 32'h3d0244a7;
8'h75 : rvCrc[25] <= 32'hdd11e7ed;
8'h76 : rvCrc[25] <= 32'hf9e41f84;
8'h77 : rvCrc[25] <= 32'h19f7bcce;
8'h78 : rvCrc[25] <= 32'haed5a503;
8'h79 : rvCrc[25] <= 32'h4ec60649;
8'h7a : rvCrc[25] <= 32'h6a33fe20;
8'h7b : rvCrc[25] <= 32'h8a205d6a;
8'h7c : rvCrc[25] <= 32'h23d80ef2;
8'h7d : rvCrc[25] <= 32'hc3cbadb8;
8'h7e : rvCrc[25] <= 32'he73e55d1;
8'h7f : rvCrc[25] <= 32'h072df69b;
8'h80 : rvCrc[25] <= 32'he965b8e7;
8'h81 : rvCrc[25] <= 32'h09761bad;
8'h82 : rvCrc[25] <= 32'h2d83e3c4;
8'h83 : rvCrc[25] <= 32'hcd90408e;
8'h84 : rvCrc[25] <= 32'h64681316;
8'h85 : rvCrc[25] <= 32'h847bb05c;
8'h86 : rvCrc[25] <= 32'ha08e4835;
8'h87 : rvCrc[25] <= 32'h409deb7f;
8'h88 : rvCrc[25] <= 32'hf7bff2b2;
8'h89 : rvCrc[25] <= 32'h17ac51f8;
8'h8a : rvCrc[25] <= 32'h3359a991;
8'h8b : rvCrc[25] <= 32'hd34a0adb;
8'h8c : rvCrc[25] <= 32'h7ab25943;
8'h8d : rvCrc[25] <= 32'h9aa1fa09;
8'h8e : rvCrc[25] <= 32'hbe540260;
8'h8f : rvCrc[25] <= 32'h5e47a12a;
8'h90 : rvCrc[25] <= 32'hd4d12c4d;
8'h91 : rvCrc[25] <= 32'h34c28f07;
8'h92 : rvCrc[25] <= 32'h1037776e;
8'h93 : rvCrc[25] <= 32'hf024d424;
8'h94 : rvCrc[25] <= 32'h59dc87bc;
8'h95 : rvCrc[25] <= 32'hb9cf24f6;
8'h96 : rvCrc[25] <= 32'h9d3adc9f;
8'h97 : rvCrc[25] <= 32'h7d297fd5;
8'h98 : rvCrc[25] <= 32'hca0b6618;
8'h99 : rvCrc[25] <= 32'h2a18c552;
8'h9a : rvCrc[25] <= 32'h0eed3d3b;
8'h9b : rvCrc[25] <= 32'heefe9e71;
8'h9c : rvCrc[25] <= 32'h4706cde9;
8'h9d : rvCrc[25] <= 32'ha7156ea3;
8'h9e : rvCrc[25] <= 32'h83e096ca;
8'h9f : rvCrc[25] <= 32'h63f33580;
8'ha0 : rvCrc[25] <= 32'h920c91b3;
8'ha1 : rvCrc[25] <= 32'h721f32f9;
8'ha2 : rvCrc[25] <= 32'h56eaca90;
8'ha3 : rvCrc[25] <= 32'hb6f969da;
8'ha4 : rvCrc[25] <= 32'h1f013a42;
8'ha5 : rvCrc[25] <= 32'hff129908;
8'ha6 : rvCrc[25] <= 32'hdbe76161;
8'ha7 : rvCrc[25] <= 32'h3bf4c22b;
8'ha8 : rvCrc[25] <= 32'h8cd6dbe6;
8'ha9 : rvCrc[25] <= 32'h6cc578ac;
8'haa : rvCrc[25] <= 32'h483080c5;
8'hab : rvCrc[25] <= 32'ha823238f;
8'hac : rvCrc[25] <= 32'h01db7017;
8'had : rvCrc[25] <= 32'he1c8d35d;
8'hae : rvCrc[25] <= 32'hc53d2b34;
8'haf : rvCrc[25] <= 32'h252e887e;
8'hb0 : rvCrc[25] <= 32'hafb80519;
8'hb1 : rvCrc[25] <= 32'h4faba653;
8'hb2 : rvCrc[25] <= 32'h6b5e5e3a;
8'hb3 : rvCrc[25] <= 32'h8b4dfd70;
8'hb4 : rvCrc[25] <= 32'h22b5aee8;
8'hb5 : rvCrc[25] <= 32'hc2a60da2;
8'hb6 : rvCrc[25] <= 32'he653f5cb;
8'hb7 : rvCrc[25] <= 32'h06405681;
8'hb8 : rvCrc[25] <= 32'hb1624f4c;
8'hb9 : rvCrc[25] <= 32'h5171ec06;
8'hba : rvCrc[25] <= 32'h7584146f;
8'hbb : rvCrc[25] <= 32'h9597b725;
8'hbc : rvCrc[25] <= 32'h3c6fe4bd;
8'hbd : rvCrc[25] <= 32'hdc7c47f7;
8'hbe : rvCrc[25] <= 32'hf889bf9e;
8'hbf : rvCrc[25] <= 32'h189a1cd4;
8'hc0 : rvCrc[25] <= 32'h1fb7ea4f;
8'hc1 : rvCrc[25] <= 32'hffa44905;
8'hc2 : rvCrc[25] <= 32'hdb51b16c;
8'hc3 : rvCrc[25] <= 32'h3b421226;
8'hc4 : rvCrc[25] <= 32'h92ba41be;
8'hc5 : rvCrc[25] <= 32'h72a9e2f4;
8'hc6 : rvCrc[25] <= 32'h565c1a9d;
8'hc7 : rvCrc[25] <= 32'hb64fb9d7;
8'hc8 : rvCrc[25] <= 32'h016da01a;
8'hc9 : rvCrc[25] <= 32'he17e0350;
8'hca : rvCrc[25] <= 32'hc58bfb39;
8'hcb : rvCrc[25] <= 32'h25985873;
8'hcc : rvCrc[25] <= 32'h8c600beb;
8'hcd : rvCrc[25] <= 32'h6c73a8a1;
8'hce : rvCrc[25] <= 32'h488650c8;
8'hcf : rvCrc[25] <= 32'ha895f382;
8'hd0 : rvCrc[25] <= 32'h22037ee5;
8'hd1 : rvCrc[25] <= 32'hc210ddaf;
8'hd2 : rvCrc[25] <= 32'he6e525c6;
8'hd3 : rvCrc[25] <= 32'h06f6868c;
8'hd4 : rvCrc[25] <= 32'haf0ed514;
8'hd5 : rvCrc[25] <= 32'h4f1d765e;
8'hd6 : rvCrc[25] <= 32'h6be88e37;
8'hd7 : rvCrc[25] <= 32'h8bfb2d7d;
8'hd8 : rvCrc[25] <= 32'h3cd934b0;
8'hd9 : rvCrc[25] <= 32'hdcca97fa;
8'hda : rvCrc[25] <= 32'hf83f6f93;
8'hdb : rvCrc[25] <= 32'h182cccd9;
8'hdc : rvCrc[25] <= 32'hb1d49f41;
8'hdd : rvCrc[25] <= 32'h51c73c0b;
8'hde : rvCrc[25] <= 32'h7532c462;
8'hdf : rvCrc[25] <= 32'h95216728;
8'he0 : rvCrc[25] <= 32'h64dec31b;
8'he1 : rvCrc[25] <= 32'h84cd6051;
8'he2 : rvCrc[25] <= 32'ha0389838;
8'he3 : rvCrc[25] <= 32'h402b3b72;
8'he4 : rvCrc[25] <= 32'he9d368ea;
8'he5 : rvCrc[25] <= 32'h09c0cba0;
8'he6 : rvCrc[25] <= 32'h2d3533c9;
8'he7 : rvCrc[25] <= 32'hcd269083;
8'he8 : rvCrc[25] <= 32'h7a04894e;
8'he9 : rvCrc[25] <= 32'h9a172a04;
8'hea : rvCrc[25] <= 32'hbee2d26d;
8'heb : rvCrc[25] <= 32'h5ef17127;
8'hec : rvCrc[25] <= 32'hf70922bf;
8'hed : rvCrc[25] <= 32'h171a81f5;
8'hee : rvCrc[25] <= 32'h33ef799c;
8'hef : rvCrc[25] <= 32'hd3fcdad6;
8'hf0 : rvCrc[25] <= 32'h596a57b1;
8'hf1 : rvCrc[25] <= 32'hb979f4fb;
8'hf2 : rvCrc[25] <= 32'h9d8c0c92;
8'hf3 : rvCrc[25] <= 32'h7d9fafd8;
8'hf4 : rvCrc[25] <= 32'hd467fc40;
8'hf5 : rvCrc[25] <= 32'h34745f0a;
8'hf6 : rvCrc[25] <= 32'h1081a763;
8'hf7 : rvCrc[25] <= 32'hf0920429;
8'hf8 : rvCrc[25] <= 32'h47b01de4;
8'hf9 : rvCrc[25] <= 32'ha7a3beae;
8'hfa : rvCrc[25] <= 32'h835646c7;
8'hfb : rvCrc[25] <= 32'h6345e58d;
8'hfc : rvCrc[25] <= 32'hcabdb615;
8'hfd : rvCrc[25] <= 32'h2aae155f;
8'hfe : rvCrc[25] <= 32'h0e5bed36;
8'hff : rvCrc[25] <= 32'hee484e7c;
endcase
case(iv_Input[215:208])
8'h00 : rvCrc[26] <= 32'h00000000;
8'h01 : rvCrc[26] <= 32'hd60a6c79;
8'h02 : rvCrc[26] <= 32'ha8d5c545;
8'h03 : rvCrc[26] <= 32'h7edfa93c;
8'h04 : rvCrc[26] <= 32'h556a973d;
8'h05 : rvCrc[26] <= 32'h8360fb44;
8'h06 : rvCrc[26] <= 32'hfdbf5278;
8'h07 : rvCrc[26] <= 32'h2bb53e01;
8'h08 : rvCrc[26] <= 32'haad52e7a;
8'h09 : rvCrc[26] <= 32'h7cdf4203;
8'h0a : rvCrc[26] <= 32'h0200eb3f;
8'h0b : rvCrc[26] <= 32'hd40a8746;
8'h0c : rvCrc[26] <= 32'hffbfb947;
8'h0d : rvCrc[26] <= 32'h29b5d53e;
8'h0e : rvCrc[26] <= 32'h576a7c02;
8'h0f : rvCrc[26] <= 32'h8160107b;
8'h10 : rvCrc[26] <= 32'h516b4143;
8'h11 : rvCrc[26] <= 32'h87612d3a;
8'h12 : rvCrc[26] <= 32'hf9be8406;
8'h13 : rvCrc[26] <= 32'h2fb4e87f;
8'h14 : rvCrc[26] <= 32'h0401d67e;
8'h15 : rvCrc[26] <= 32'hd20bba07;
8'h16 : rvCrc[26] <= 32'hacd4133b;
8'h17 : rvCrc[26] <= 32'h7ade7f42;
8'h18 : rvCrc[26] <= 32'hfbbe6f39;
8'h19 : rvCrc[26] <= 32'h2db40340;
8'h1a : rvCrc[26] <= 32'h536baa7c;
8'h1b : rvCrc[26] <= 32'h8561c605;
8'h1c : rvCrc[26] <= 32'haed4f804;
8'h1d : rvCrc[26] <= 32'h78de947d;
8'h1e : rvCrc[26] <= 32'h06013d41;
8'h1f : rvCrc[26] <= 32'hd00b5138;
8'h20 : rvCrc[26] <= 32'ha2d68286;
8'h21 : rvCrc[26] <= 32'h74dceeff;
8'h22 : rvCrc[26] <= 32'h0a0347c3;
8'h23 : rvCrc[26] <= 32'hdc092bba;
8'h24 : rvCrc[26] <= 32'hf7bc15bb;
8'h25 : rvCrc[26] <= 32'h21b679c2;
8'h26 : rvCrc[26] <= 32'h5f69d0fe;
8'h27 : rvCrc[26] <= 32'h8963bc87;
8'h28 : rvCrc[26] <= 32'h0803acfc;
8'h29 : rvCrc[26] <= 32'hde09c085;
8'h2a : rvCrc[26] <= 32'ha0d669b9;
8'h2b : rvCrc[26] <= 32'h76dc05c0;
8'h2c : rvCrc[26] <= 32'h5d693bc1;
8'h2d : rvCrc[26] <= 32'h8b6357b8;
8'h2e : rvCrc[26] <= 32'hf5bcfe84;
8'h2f : rvCrc[26] <= 32'h23b692fd;
8'h30 : rvCrc[26] <= 32'hf3bdc3c5;
8'h31 : rvCrc[26] <= 32'h25b7afbc;
8'h32 : rvCrc[26] <= 32'h5b680680;
8'h33 : rvCrc[26] <= 32'h8d626af9;
8'h34 : rvCrc[26] <= 32'ha6d754f8;
8'h35 : rvCrc[26] <= 32'h70dd3881;
8'h36 : rvCrc[26] <= 32'h0e0291bd;
8'h37 : rvCrc[26] <= 32'hd808fdc4;
8'h38 : rvCrc[26] <= 32'h5968edbf;
8'h39 : rvCrc[26] <= 32'h8f6281c6;
8'h3a : rvCrc[26] <= 32'hf1bd28fa;
8'h3b : rvCrc[26] <= 32'h27b74483;
8'h3c : rvCrc[26] <= 32'h0c027a82;
8'h3d : rvCrc[26] <= 32'hda0816fb;
8'h3e : rvCrc[26] <= 32'ha4d7bfc7;
8'h3f : rvCrc[26] <= 32'h72ddd3be;
8'h40 : rvCrc[26] <= 32'h416c18bb;
8'h41 : rvCrc[26] <= 32'h976674c2;
8'h42 : rvCrc[26] <= 32'he9b9ddfe;
8'h43 : rvCrc[26] <= 32'h3fb3b187;
8'h44 : rvCrc[26] <= 32'h14068f86;
8'h45 : rvCrc[26] <= 32'hc20ce3ff;
8'h46 : rvCrc[26] <= 32'hbcd34ac3;
8'h47 : rvCrc[26] <= 32'h6ad926ba;
8'h48 : rvCrc[26] <= 32'hebb936c1;
8'h49 : rvCrc[26] <= 32'h3db35ab8;
8'h4a : rvCrc[26] <= 32'h436cf384;
8'h4b : rvCrc[26] <= 32'h95669ffd;
8'h4c : rvCrc[26] <= 32'hbed3a1fc;
8'h4d : rvCrc[26] <= 32'h68d9cd85;
8'h4e : rvCrc[26] <= 32'h160664b9;
8'h4f : rvCrc[26] <= 32'hc00c08c0;
8'h50 : rvCrc[26] <= 32'h100759f8;
8'h51 : rvCrc[26] <= 32'hc60d3581;
8'h52 : rvCrc[26] <= 32'hb8d29cbd;
8'h53 : rvCrc[26] <= 32'h6ed8f0c4;
8'h54 : rvCrc[26] <= 32'h456dcec5;
8'h55 : rvCrc[26] <= 32'h9367a2bc;
8'h56 : rvCrc[26] <= 32'hedb80b80;
8'h57 : rvCrc[26] <= 32'h3bb267f9;
8'h58 : rvCrc[26] <= 32'hbad27782;
8'h59 : rvCrc[26] <= 32'h6cd81bfb;
8'h5a : rvCrc[26] <= 32'h1207b2c7;
8'h5b : rvCrc[26] <= 32'hc40ddebe;
8'h5c : rvCrc[26] <= 32'hefb8e0bf;
8'h5d : rvCrc[26] <= 32'h39b28cc6;
8'h5e : rvCrc[26] <= 32'h476d25fa;
8'h5f : rvCrc[26] <= 32'h91674983;
8'h60 : rvCrc[26] <= 32'he3ba9a3d;
8'h61 : rvCrc[26] <= 32'h35b0f644;
8'h62 : rvCrc[26] <= 32'h4b6f5f78;
8'h63 : rvCrc[26] <= 32'h9d653301;
8'h64 : rvCrc[26] <= 32'hb6d00d00;
8'h65 : rvCrc[26] <= 32'h60da6179;
8'h66 : rvCrc[26] <= 32'h1e05c845;
8'h67 : rvCrc[26] <= 32'hc80fa43c;
8'h68 : rvCrc[26] <= 32'h496fb447;
8'h69 : rvCrc[26] <= 32'h9f65d83e;
8'h6a : rvCrc[26] <= 32'he1ba7102;
8'h6b : rvCrc[26] <= 32'h37b01d7b;
8'h6c : rvCrc[26] <= 32'h1c05237a;
8'h6d : rvCrc[26] <= 32'hca0f4f03;
8'h6e : rvCrc[26] <= 32'hb4d0e63f;
8'h6f : rvCrc[26] <= 32'h62da8a46;
8'h70 : rvCrc[26] <= 32'hb2d1db7e;
8'h71 : rvCrc[26] <= 32'h64dbb707;
8'h72 : rvCrc[26] <= 32'h1a041e3b;
8'h73 : rvCrc[26] <= 32'hcc0e7242;
8'h74 : rvCrc[26] <= 32'he7bb4c43;
8'h75 : rvCrc[26] <= 32'h31b1203a;
8'h76 : rvCrc[26] <= 32'h4f6e8906;
8'h77 : rvCrc[26] <= 32'h9964e57f;
8'h78 : rvCrc[26] <= 32'h1804f504;
8'h79 : rvCrc[26] <= 32'hce0e997d;
8'h7a : rvCrc[26] <= 32'hb0d13041;
8'h7b : rvCrc[26] <= 32'h66db5c38;
8'h7c : rvCrc[26] <= 32'h4d6e6239;
8'h7d : rvCrc[26] <= 32'h9b640e40;
8'h7e : rvCrc[26] <= 32'he5bba77c;
8'h7f : rvCrc[26] <= 32'h33b1cb05;
8'h80 : rvCrc[26] <= 32'h82d83176;
8'h81 : rvCrc[26] <= 32'h54d25d0f;
8'h82 : rvCrc[26] <= 32'h2a0df433;
8'h83 : rvCrc[26] <= 32'hfc07984a;
8'h84 : rvCrc[26] <= 32'hd7b2a64b;
8'h85 : rvCrc[26] <= 32'h01b8ca32;
8'h86 : rvCrc[26] <= 32'h7f67630e;
8'h87 : rvCrc[26] <= 32'ha96d0f77;
8'h88 : rvCrc[26] <= 32'h280d1f0c;
8'h89 : rvCrc[26] <= 32'hfe077375;
8'h8a : rvCrc[26] <= 32'h80d8da49;
8'h8b : rvCrc[26] <= 32'h56d2b630;
8'h8c : rvCrc[26] <= 32'h7d678831;
8'h8d : rvCrc[26] <= 32'hab6de448;
8'h8e : rvCrc[26] <= 32'hd5b24d74;
8'h8f : rvCrc[26] <= 32'h03b8210d;
8'h90 : rvCrc[26] <= 32'hd3b37035;
8'h91 : rvCrc[26] <= 32'h05b91c4c;
8'h92 : rvCrc[26] <= 32'h7b66b570;
8'h93 : rvCrc[26] <= 32'had6cd909;
8'h94 : rvCrc[26] <= 32'h86d9e708;
8'h95 : rvCrc[26] <= 32'h50d38b71;
8'h96 : rvCrc[26] <= 32'h2e0c224d;
8'h97 : rvCrc[26] <= 32'hf8064e34;
8'h98 : rvCrc[26] <= 32'h79665e4f;
8'h99 : rvCrc[26] <= 32'haf6c3236;
8'h9a : rvCrc[26] <= 32'hd1b39b0a;
8'h9b : rvCrc[26] <= 32'h07b9f773;
8'h9c : rvCrc[26] <= 32'h2c0cc972;
8'h9d : rvCrc[26] <= 32'hfa06a50b;
8'h9e : rvCrc[26] <= 32'h84d90c37;
8'h9f : rvCrc[26] <= 32'h52d3604e;
8'ha0 : rvCrc[26] <= 32'h200eb3f0;
8'ha1 : rvCrc[26] <= 32'hf604df89;
8'ha2 : rvCrc[26] <= 32'h88db76b5;
8'ha3 : rvCrc[26] <= 32'h5ed11acc;
8'ha4 : rvCrc[26] <= 32'h756424cd;
8'ha5 : rvCrc[26] <= 32'ha36e48b4;
8'ha6 : rvCrc[26] <= 32'hddb1e188;
8'ha7 : rvCrc[26] <= 32'h0bbb8df1;
8'ha8 : rvCrc[26] <= 32'h8adb9d8a;
8'ha9 : rvCrc[26] <= 32'h5cd1f1f3;
8'haa : rvCrc[26] <= 32'h220e58cf;
8'hab : rvCrc[26] <= 32'hf40434b6;
8'hac : rvCrc[26] <= 32'hdfb10ab7;
8'had : rvCrc[26] <= 32'h09bb66ce;
8'hae : rvCrc[26] <= 32'h7764cff2;
8'haf : rvCrc[26] <= 32'ha16ea38b;
8'hb0 : rvCrc[26] <= 32'h7165f2b3;
8'hb1 : rvCrc[26] <= 32'ha76f9eca;
8'hb2 : rvCrc[26] <= 32'hd9b037f6;
8'hb3 : rvCrc[26] <= 32'h0fba5b8f;
8'hb4 : rvCrc[26] <= 32'h240f658e;
8'hb5 : rvCrc[26] <= 32'hf20509f7;
8'hb6 : rvCrc[26] <= 32'h8cdaa0cb;
8'hb7 : rvCrc[26] <= 32'h5ad0ccb2;
8'hb8 : rvCrc[26] <= 32'hdbb0dcc9;
8'hb9 : rvCrc[26] <= 32'h0dbab0b0;
8'hba : rvCrc[26] <= 32'h7365198c;
8'hbb : rvCrc[26] <= 32'ha56f75f5;
8'hbc : rvCrc[26] <= 32'h8eda4bf4;
8'hbd : rvCrc[26] <= 32'h58d0278d;
8'hbe : rvCrc[26] <= 32'h260f8eb1;
8'hbf : rvCrc[26] <= 32'hf005e2c8;
8'hc0 : rvCrc[26] <= 32'hc3b429cd;
8'hc1 : rvCrc[26] <= 32'h15be45b4;
8'hc2 : rvCrc[26] <= 32'h6b61ec88;
8'hc3 : rvCrc[26] <= 32'hbd6b80f1;
8'hc4 : rvCrc[26] <= 32'h96debef0;
8'hc5 : rvCrc[26] <= 32'h40d4d289;
8'hc6 : rvCrc[26] <= 32'h3e0b7bb5;
8'hc7 : rvCrc[26] <= 32'he80117cc;
8'hc8 : rvCrc[26] <= 32'h696107b7;
8'hc9 : rvCrc[26] <= 32'hbf6b6bce;
8'hca : rvCrc[26] <= 32'hc1b4c2f2;
8'hcb : rvCrc[26] <= 32'h17beae8b;
8'hcc : rvCrc[26] <= 32'h3c0b908a;
8'hcd : rvCrc[26] <= 32'hea01fcf3;
8'hce : rvCrc[26] <= 32'h94de55cf;
8'hcf : rvCrc[26] <= 32'h42d439b6;
8'hd0 : rvCrc[26] <= 32'h92df688e;
8'hd1 : rvCrc[26] <= 32'h44d504f7;
8'hd2 : rvCrc[26] <= 32'h3a0aadcb;
8'hd3 : rvCrc[26] <= 32'hec00c1b2;
8'hd4 : rvCrc[26] <= 32'hc7b5ffb3;
8'hd5 : rvCrc[26] <= 32'h11bf93ca;
8'hd6 : rvCrc[26] <= 32'h6f603af6;
8'hd7 : rvCrc[26] <= 32'hb96a568f;
8'hd8 : rvCrc[26] <= 32'h380a46f4;
8'hd9 : rvCrc[26] <= 32'hee002a8d;
8'hda : rvCrc[26] <= 32'h90df83b1;
8'hdb : rvCrc[26] <= 32'h46d5efc8;
8'hdc : rvCrc[26] <= 32'h6d60d1c9;
8'hdd : rvCrc[26] <= 32'hbb6abdb0;
8'hde : rvCrc[26] <= 32'hc5b5148c;
8'hdf : rvCrc[26] <= 32'h13bf78f5;
8'he0 : rvCrc[26] <= 32'h6162ab4b;
8'he1 : rvCrc[26] <= 32'hb768c732;
8'he2 : rvCrc[26] <= 32'hc9b76e0e;
8'he3 : rvCrc[26] <= 32'h1fbd0277;
8'he4 : rvCrc[26] <= 32'h34083c76;
8'he5 : rvCrc[26] <= 32'he202500f;
8'he6 : rvCrc[26] <= 32'h9cddf933;
8'he7 : rvCrc[26] <= 32'h4ad7954a;
8'he8 : rvCrc[26] <= 32'hcbb78531;
8'he9 : rvCrc[26] <= 32'h1dbde948;
8'hea : rvCrc[26] <= 32'h63624074;
8'heb : rvCrc[26] <= 32'hb5682c0d;
8'hec : rvCrc[26] <= 32'h9edd120c;
8'hed : rvCrc[26] <= 32'h48d77e75;
8'hee : rvCrc[26] <= 32'h3608d749;
8'hef : rvCrc[26] <= 32'he002bb30;
8'hf0 : rvCrc[26] <= 32'h3009ea08;
8'hf1 : rvCrc[26] <= 32'he6038671;
8'hf2 : rvCrc[26] <= 32'h98dc2f4d;
8'hf3 : rvCrc[26] <= 32'h4ed64334;
8'hf4 : rvCrc[26] <= 32'h65637d35;
8'hf5 : rvCrc[26] <= 32'hb369114c;
8'hf6 : rvCrc[26] <= 32'hcdb6b870;
8'hf7 : rvCrc[26] <= 32'h1bbcd409;
8'hf8 : rvCrc[26] <= 32'h9adcc472;
8'hf9 : rvCrc[26] <= 32'h4cd6a80b;
8'hfa : rvCrc[26] <= 32'h32090137;
8'hfb : rvCrc[26] <= 32'he4036d4e;
8'hfc : rvCrc[26] <= 32'hcfb6534f;
8'hfd : rvCrc[26] <= 32'h19bc3f36;
8'hfe : rvCrc[26] <= 32'h6763960a;
8'hff : rvCrc[26] <= 32'hb169fa73;
endcase
case(iv_Input[223:216])
8'h00 : rvCrc[27] <= 32'h00000000;
8'h01 : rvCrc[27] <= 32'h01717f5b;
8'h02 : rvCrc[27] <= 32'h02e2feb6;
8'h03 : rvCrc[27] <= 32'h039381ed;
8'h04 : rvCrc[27] <= 32'h05c5fd6c;
8'h05 : rvCrc[27] <= 32'h04b48237;
8'h06 : rvCrc[27] <= 32'h072703da;
8'h07 : rvCrc[27] <= 32'h06567c81;
8'h08 : rvCrc[27] <= 32'h0b8bfad8;
8'h09 : rvCrc[27] <= 32'h0afa8583;
8'h0a : rvCrc[27] <= 32'h0969046e;
8'h0b : rvCrc[27] <= 32'h08187b35;
8'h0c : rvCrc[27] <= 32'h0e4e07b4;
8'h0d : rvCrc[27] <= 32'h0f3f78ef;
8'h0e : rvCrc[27] <= 32'h0cacf902;
8'h0f : rvCrc[27] <= 32'h0ddd8659;
8'h10 : rvCrc[27] <= 32'h1717f5b0;
8'h11 : rvCrc[27] <= 32'h16668aeb;
8'h12 : rvCrc[27] <= 32'h15f50b06;
8'h13 : rvCrc[27] <= 32'h1484745d;
8'h14 : rvCrc[27] <= 32'h12d208dc;
8'h15 : rvCrc[27] <= 32'h13a37787;
8'h16 : rvCrc[27] <= 32'h1030f66a;
8'h17 : rvCrc[27] <= 32'h11418931;
8'h18 : rvCrc[27] <= 32'h1c9c0f68;
8'h19 : rvCrc[27] <= 32'h1ded7033;
8'h1a : rvCrc[27] <= 32'h1e7ef1de;
8'h1b : rvCrc[27] <= 32'h1f0f8e85;
8'h1c : rvCrc[27] <= 32'h1959f204;
8'h1d : rvCrc[27] <= 32'h18288d5f;
8'h1e : rvCrc[27] <= 32'h1bbb0cb2;
8'h1f : rvCrc[27] <= 32'h1aca73e9;
8'h20 : rvCrc[27] <= 32'h2e2feb60;
8'h21 : rvCrc[27] <= 32'h2f5e943b;
8'h22 : rvCrc[27] <= 32'h2ccd15d6;
8'h23 : rvCrc[27] <= 32'h2dbc6a8d;
8'h24 : rvCrc[27] <= 32'h2bea160c;
8'h25 : rvCrc[27] <= 32'h2a9b6957;
8'h26 : rvCrc[27] <= 32'h2908e8ba;
8'h27 : rvCrc[27] <= 32'h287997e1;
8'h28 : rvCrc[27] <= 32'h25a411b8;
8'h29 : rvCrc[27] <= 32'h24d56ee3;
8'h2a : rvCrc[27] <= 32'h2746ef0e;
8'h2b : rvCrc[27] <= 32'h26379055;
8'h2c : rvCrc[27] <= 32'h2061ecd4;
8'h2d : rvCrc[27] <= 32'h2110938f;
8'h2e : rvCrc[27] <= 32'h22831262;
8'h2f : rvCrc[27] <= 32'h23f26d39;
8'h30 : rvCrc[27] <= 32'h39381ed0;
8'h31 : rvCrc[27] <= 32'h3849618b;
8'h32 : rvCrc[27] <= 32'h3bdae066;
8'h33 : rvCrc[27] <= 32'h3aab9f3d;
8'h34 : rvCrc[27] <= 32'h3cfde3bc;
8'h35 : rvCrc[27] <= 32'h3d8c9ce7;
8'h36 : rvCrc[27] <= 32'h3e1f1d0a;
8'h37 : rvCrc[27] <= 32'h3f6e6251;
8'h38 : rvCrc[27] <= 32'h32b3e408;
8'h39 : rvCrc[27] <= 32'h33c29b53;
8'h3a : rvCrc[27] <= 32'h30511abe;
8'h3b : rvCrc[27] <= 32'h312065e5;
8'h3c : rvCrc[27] <= 32'h37761964;
8'h3d : rvCrc[27] <= 32'h3607663f;
8'h3e : rvCrc[27] <= 32'h3594e7d2;
8'h3f : rvCrc[27] <= 32'h34e59889;
8'h40 : rvCrc[27] <= 32'h5c5fd6c0;
8'h41 : rvCrc[27] <= 32'h5d2ea99b;
8'h42 : rvCrc[27] <= 32'h5ebd2876;
8'h43 : rvCrc[27] <= 32'h5fcc572d;
8'h44 : rvCrc[27] <= 32'h599a2bac;
8'h45 : rvCrc[27] <= 32'h58eb54f7;
8'h46 : rvCrc[27] <= 32'h5b78d51a;
8'h47 : rvCrc[27] <= 32'h5a09aa41;
8'h48 : rvCrc[27] <= 32'h57d42c18;
8'h49 : rvCrc[27] <= 32'h56a55343;
8'h4a : rvCrc[27] <= 32'h5536d2ae;
8'h4b : rvCrc[27] <= 32'h5447adf5;
8'h4c : rvCrc[27] <= 32'h5211d174;
8'h4d : rvCrc[27] <= 32'h5360ae2f;
8'h4e : rvCrc[27] <= 32'h50f32fc2;
8'h4f : rvCrc[27] <= 32'h51825099;
8'h50 : rvCrc[27] <= 32'h4b482370;
8'h51 : rvCrc[27] <= 32'h4a395c2b;
8'h52 : rvCrc[27] <= 32'h49aaddc6;
8'h53 : rvCrc[27] <= 32'h48dba29d;
8'h54 : rvCrc[27] <= 32'h4e8dde1c;
8'h55 : rvCrc[27] <= 32'h4ffca147;
8'h56 : rvCrc[27] <= 32'h4c6f20aa;
8'h57 : rvCrc[27] <= 32'h4d1e5ff1;
8'h58 : rvCrc[27] <= 32'h40c3d9a8;
8'h59 : rvCrc[27] <= 32'h41b2a6f3;
8'h5a : rvCrc[27] <= 32'h4221271e;
8'h5b : rvCrc[27] <= 32'h43505845;
8'h5c : rvCrc[27] <= 32'h450624c4;
8'h5d : rvCrc[27] <= 32'h44775b9f;
8'h5e : rvCrc[27] <= 32'h47e4da72;
8'h5f : rvCrc[27] <= 32'h4695a529;
8'h60 : rvCrc[27] <= 32'h72703da0;
8'h61 : rvCrc[27] <= 32'h730142fb;
8'h62 : rvCrc[27] <= 32'h7092c316;
8'h63 : rvCrc[27] <= 32'h71e3bc4d;
8'h64 : rvCrc[27] <= 32'h77b5c0cc;
8'h65 : rvCrc[27] <= 32'h76c4bf97;
8'h66 : rvCrc[27] <= 32'h75573e7a;
8'h67 : rvCrc[27] <= 32'h74264121;
8'h68 : rvCrc[27] <= 32'h79fbc778;
8'h69 : rvCrc[27] <= 32'h788ab823;
8'h6a : rvCrc[27] <= 32'h7b1939ce;
8'h6b : rvCrc[27] <= 32'h7a684695;
8'h6c : rvCrc[27] <= 32'h7c3e3a14;
8'h6d : rvCrc[27] <= 32'h7d4f454f;
8'h6e : rvCrc[27] <= 32'h7edcc4a2;
8'h6f : rvCrc[27] <= 32'h7fadbbf9;
8'h70 : rvCrc[27] <= 32'h6567c810;
8'h71 : rvCrc[27] <= 32'h6416b74b;
8'h72 : rvCrc[27] <= 32'h678536a6;
8'h73 : rvCrc[27] <= 32'h66f449fd;
8'h74 : rvCrc[27] <= 32'h60a2357c;
8'h75 : rvCrc[27] <= 32'h61d34a27;
8'h76 : rvCrc[27] <= 32'h6240cbca;
8'h77 : rvCrc[27] <= 32'h6331b491;
8'h78 : rvCrc[27] <= 32'h6eec32c8;
8'h79 : rvCrc[27] <= 32'h6f9d4d93;
8'h7a : rvCrc[27] <= 32'h6c0ecc7e;
8'h7b : rvCrc[27] <= 32'h6d7fb325;
8'h7c : rvCrc[27] <= 32'h6b29cfa4;
8'h7d : rvCrc[27] <= 32'h6a58b0ff;
8'h7e : rvCrc[27] <= 32'h69cb3112;
8'h7f : rvCrc[27] <= 32'h68ba4e49;
8'h80 : rvCrc[27] <= 32'hb8bfad80;
8'h81 : rvCrc[27] <= 32'hb9ced2db;
8'h82 : rvCrc[27] <= 32'hba5d5336;
8'h83 : rvCrc[27] <= 32'hbb2c2c6d;
8'h84 : rvCrc[27] <= 32'hbd7a50ec;
8'h85 : rvCrc[27] <= 32'hbc0b2fb7;
8'h86 : rvCrc[27] <= 32'hbf98ae5a;
8'h87 : rvCrc[27] <= 32'hbee9d101;
8'h88 : rvCrc[27] <= 32'hb3345758;
8'h89 : rvCrc[27] <= 32'hb2452803;
8'h8a : rvCrc[27] <= 32'hb1d6a9ee;
8'h8b : rvCrc[27] <= 32'hb0a7d6b5;
8'h8c : rvCrc[27] <= 32'hb6f1aa34;
8'h8d : rvCrc[27] <= 32'hb780d56f;
8'h8e : rvCrc[27] <= 32'hb4135482;
8'h8f : rvCrc[27] <= 32'hb5622bd9;
8'h90 : rvCrc[27] <= 32'hafa85830;
8'h91 : rvCrc[27] <= 32'haed9276b;
8'h92 : rvCrc[27] <= 32'had4aa686;
8'h93 : rvCrc[27] <= 32'hac3bd9dd;
8'h94 : rvCrc[27] <= 32'haa6da55c;
8'h95 : rvCrc[27] <= 32'hab1cda07;
8'h96 : rvCrc[27] <= 32'ha88f5bea;
8'h97 : rvCrc[27] <= 32'ha9fe24b1;
8'h98 : rvCrc[27] <= 32'ha423a2e8;
8'h99 : rvCrc[27] <= 32'ha552ddb3;
8'h9a : rvCrc[27] <= 32'ha6c15c5e;
8'h9b : rvCrc[27] <= 32'ha7b02305;
8'h9c : rvCrc[27] <= 32'ha1e65f84;
8'h9d : rvCrc[27] <= 32'ha09720df;
8'h9e : rvCrc[27] <= 32'ha304a132;
8'h9f : rvCrc[27] <= 32'ha275de69;
8'ha0 : rvCrc[27] <= 32'h969046e0;
8'ha1 : rvCrc[27] <= 32'h97e139bb;
8'ha2 : rvCrc[27] <= 32'h9472b856;
8'ha3 : rvCrc[27] <= 32'h9503c70d;
8'ha4 : rvCrc[27] <= 32'h9355bb8c;
8'ha5 : rvCrc[27] <= 32'h9224c4d7;
8'ha6 : rvCrc[27] <= 32'h91b7453a;
8'ha7 : rvCrc[27] <= 32'h90c63a61;
8'ha8 : rvCrc[27] <= 32'h9d1bbc38;
8'ha9 : rvCrc[27] <= 32'h9c6ac363;
8'haa : rvCrc[27] <= 32'h9ff9428e;
8'hab : rvCrc[27] <= 32'h9e883dd5;
8'hac : rvCrc[27] <= 32'h98de4154;
8'had : rvCrc[27] <= 32'h99af3e0f;
8'hae : rvCrc[27] <= 32'h9a3cbfe2;
8'haf : rvCrc[27] <= 32'h9b4dc0b9;
8'hb0 : rvCrc[27] <= 32'h8187b350;
8'hb1 : rvCrc[27] <= 32'h80f6cc0b;
8'hb2 : rvCrc[27] <= 32'h83654de6;
8'hb3 : rvCrc[27] <= 32'h821432bd;
8'hb4 : rvCrc[27] <= 32'h84424e3c;
8'hb5 : rvCrc[27] <= 32'h85333167;
8'hb6 : rvCrc[27] <= 32'h86a0b08a;
8'hb7 : rvCrc[27] <= 32'h87d1cfd1;
8'hb8 : rvCrc[27] <= 32'h8a0c4988;
8'hb9 : rvCrc[27] <= 32'h8b7d36d3;
8'hba : rvCrc[27] <= 32'h88eeb73e;
8'hbb : rvCrc[27] <= 32'h899fc865;
8'hbc : rvCrc[27] <= 32'h8fc9b4e4;
8'hbd : rvCrc[27] <= 32'h8eb8cbbf;
8'hbe : rvCrc[27] <= 32'h8d2b4a52;
8'hbf : rvCrc[27] <= 32'h8c5a3509;
8'hc0 : rvCrc[27] <= 32'he4e07b40;
8'hc1 : rvCrc[27] <= 32'he591041b;
8'hc2 : rvCrc[27] <= 32'he60285f6;
8'hc3 : rvCrc[27] <= 32'he773faad;
8'hc4 : rvCrc[27] <= 32'he125862c;
8'hc5 : rvCrc[27] <= 32'he054f977;
8'hc6 : rvCrc[27] <= 32'he3c7789a;
8'hc7 : rvCrc[27] <= 32'he2b607c1;
8'hc8 : rvCrc[27] <= 32'hef6b8198;
8'hc9 : rvCrc[27] <= 32'hee1afec3;
8'hca : rvCrc[27] <= 32'hed897f2e;
8'hcb : rvCrc[27] <= 32'hecf80075;
8'hcc : rvCrc[27] <= 32'heaae7cf4;
8'hcd : rvCrc[27] <= 32'hebdf03af;
8'hce : rvCrc[27] <= 32'he84c8242;
8'hcf : rvCrc[27] <= 32'he93dfd19;
8'hd0 : rvCrc[27] <= 32'hf3f78ef0;
8'hd1 : rvCrc[27] <= 32'hf286f1ab;
8'hd2 : rvCrc[27] <= 32'hf1157046;
8'hd3 : rvCrc[27] <= 32'hf0640f1d;
8'hd4 : rvCrc[27] <= 32'hf632739c;
8'hd5 : rvCrc[27] <= 32'hf7430cc7;
8'hd6 : rvCrc[27] <= 32'hf4d08d2a;
8'hd7 : rvCrc[27] <= 32'hf5a1f271;
8'hd8 : rvCrc[27] <= 32'hf87c7428;
8'hd9 : rvCrc[27] <= 32'hf90d0b73;
8'hda : rvCrc[27] <= 32'hfa9e8a9e;
8'hdb : rvCrc[27] <= 32'hfbeff5c5;
8'hdc : rvCrc[27] <= 32'hfdb98944;
8'hdd : rvCrc[27] <= 32'hfcc8f61f;
8'hde : rvCrc[27] <= 32'hff5b77f2;
8'hdf : rvCrc[27] <= 32'hfe2a08a9;
8'he0 : rvCrc[27] <= 32'hcacf9020;
8'he1 : rvCrc[27] <= 32'hcbbeef7b;
8'he2 : rvCrc[27] <= 32'hc82d6e96;
8'he3 : rvCrc[27] <= 32'hc95c11cd;
8'he4 : rvCrc[27] <= 32'hcf0a6d4c;
8'he5 : rvCrc[27] <= 32'hce7b1217;
8'he6 : rvCrc[27] <= 32'hcde893fa;
8'he7 : rvCrc[27] <= 32'hcc99eca1;
8'he8 : rvCrc[27] <= 32'hc1446af8;
8'he9 : rvCrc[27] <= 32'hc03515a3;
8'hea : rvCrc[27] <= 32'hc3a6944e;
8'heb : rvCrc[27] <= 32'hc2d7eb15;
8'hec : rvCrc[27] <= 32'hc4819794;
8'hed : rvCrc[27] <= 32'hc5f0e8cf;
8'hee : rvCrc[27] <= 32'hc6636922;
8'hef : rvCrc[27] <= 32'hc7121679;
8'hf0 : rvCrc[27] <= 32'hddd86590;
8'hf1 : rvCrc[27] <= 32'hdca91acb;
8'hf2 : rvCrc[27] <= 32'hdf3a9b26;
8'hf3 : rvCrc[27] <= 32'hde4be47d;
8'hf4 : rvCrc[27] <= 32'hd81d98fc;
8'hf5 : rvCrc[27] <= 32'hd96ce7a7;
8'hf6 : rvCrc[27] <= 32'hdaff664a;
8'hf7 : rvCrc[27] <= 32'hdb8e1911;
8'hf8 : rvCrc[27] <= 32'hd6539f48;
8'hf9 : rvCrc[27] <= 32'hd722e013;
8'hfa : rvCrc[27] <= 32'hd4b161fe;
8'hfb : rvCrc[27] <= 32'hd5c01ea5;
8'hfc : rvCrc[27] <= 32'hd3966224;
8'hfd : rvCrc[27] <= 32'hd2e71d7f;
8'hfe : rvCrc[27] <= 32'hd1749c92;
8'hff : rvCrc[27] <= 32'hd005e3c9;
endcase
case(iv_Input[231:224])
8'h00 : rvCrc[28] <= 32'h00000000;
8'h01 : rvCrc[28] <= 32'h75be46b7;
8'h02 : rvCrc[28] <= 32'heb7c8d6e;
8'h03 : rvCrc[28] <= 32'h9ec2cbd9;
8'h04 : rvCrc[28] <= 32'hd238076b;
8'h05 : rvCrc[28] <= 32'ha78641dc;
8'h06 : rvCrc[28] <= 32'h39448a05;
8'h07 : rvCrc[28] <= 32'h4cfaccb2;
8'h08 : rvCrc[28] <= 32'ha0b11361;
8'h09 : rvCrc[28] <= 32'hd50f55d6;
8'h0a : rvCrc[28] <= 32'h4bcd9e0f;
8'h0b : rvCrc[28] <= 32'h3e73d8b8;
8'h0c : rvCrc[28] <= 32'h7289140a;
8'h0d : rvCrc[28] <= 32'h073752bd;
8'h0e : rvCrc[28] <= 32'h99f59964;
8'h0f : rvCrc[28] <= 32'hec4bdfd3;
8'h10 : rvCrc[28] <= 32'h45a33b75;
8'h11 : rvCrc[28] <= 32'h301d7dc2;
8'h12 : rvCrc[28] <= 32'haedfb61b;
8'h13 : rvCrc[28] <= 32'hdb61f0ac;
8'h14 : rvCrc[28] <= 32'h979b3c1e;
8'h15 : rvCrc[28] <= 32'he2257aa9;
8'h16 : rvCrc[28] <= 32'h7ce7b170;
8'h17 : rvCrc[28] <= 32'h0959f7c7;
8'h18 : rvCrc[28] <= 32'he5122814;
8'h19 : rvCrc[28] <= 32'h90ac6ea3;
8'h1a : rvCrc[28] <= 32'h0e6ea57a;
8'h1b : rvCrc[28] <= 32'h7bd0e3cd;
8'h1c : rvCrc[28] <= 32'h372a2f7f;
8'h1d : rvCrc[28] <= 32'h429469c8;
8'h1e : rvCrc[28] <= 32'hdc56a211;
8'h1f : rvCrc[28] <= 32'ha9e8e4a6;
8'h20 : rvCrc[28] <= 32'h8b4676ea;
8'h21 : rvCrc[28] <= 32'hfef8305d;
8'h22 : rvCrc[28] <= 32'h603afb84;
8'h23 : rvCrc[28] <= 32'h1584bd33;
8'h24 : rvCrc[28] <= 32'h597e7181;
8'h25 : rvCrc[28] <= 32'h2cc03736;
8'h26 : rvCrc[28] <= 32'hb202fcef;
8'h27 : rvCrc[28] <= 32'hc7bcba58;
8'h28 : rvCrc[28] <= 32'h2bf7658b;
8'h29 : rvCrc[28] <= 32'h5e49233c;
8'h2a : rvCrc[28] <= 32'hc08be8e5;
8'h2b : rvCrc[28] <= 32'hb535ae52;
8'h2c : rvCrc[28] <= 32'hf9cf62e0;
8'h2d : rvCrc[28] <= 32'h8c712457;
8'h2e : rvCrc[28] <= 32'h12b3ef8e;
8'h2f : rvCrc[28] <= 32'h670da939;
8'h30 : rvCrc[28] <= 32'hcee54d9f;
8'h31 : rvCrc[28] <= 32'hbb5b0b28;
8'h32 : rvCrc[28] <= 32'h2599c0f1;
8'h33 : rvCrc[28] <= 32'h50278646;
8'h34 : rvCrc[28] <= 32'h1cdd4af4;
8'h35 : rvCrc[28] <= 32'h69630c43;
8'h36 : rvCrc[28] <= 32'hf7a1c79a;
8'h37 : rvCrc[28] <= 32'h821f812d;
8'h38 : rvCrc[28] <= 32'h6e545efe;
8'h39 : rvCrc[28] <= 32'h1bea1849;
8'h3a : rvCrc[28] <= 32'h8528d390;
8'h3b : rvCrc[28] <= 32'hf0969527;
8'h3c : rvCrc[28] <= 32'hbc6c5995;
8'h3d : rvCrc[28] <= 32'hc9d21f22;
8'h3e : rvCrc[28] <= 32'h5710d4fb;
8'h3f : rvCrc[28] <= 32'h22ae924c;
8'h40 : rvCrc[28] <= 32'h124df063;
8'h41 : rvCrc[28] <= 32'h67f3b6d4;
8'h42 : rvCrc[28] <= 32'hf9317d0d;
8'h43 : rvCrc[28] <= 32'h8c8f3bba;
8'h44 : rvCrc[28] <= 32'hc075f708;
8'h45 : rvCrc[28] <= 32'hb5cbb1bf;
8'h46 : rvCrc[28] <= 32'h2b097a66;
8'h47 : rvCrc[28] <= 32'h5eb73cd1;
8'h48 : rvCrc[28] <= 32'hb2fce302;
8'h49 : rvCrc[28] <= 32'hc742a5b5;
8'h4a : rvCrc[28] <= 32'h59806e6c;
8'h4b : rvCrc[28] <= 32'h2c3e28db;
8'h4c : rvCrc[28] <= 32'h60c4e469;
8'h4d : rvCrc[28] <= 32'h157aa2de;
8'h4e : rvCrc[28] <= 32'h8bb86907;
8'h4f : rvCrc[28] <= 32'hfe062fb0;
8'h50 : rvCrc[28] <= 32'h57eecb16;
8'h51 : rvCrc[28] <= 32'h22508da1;
8'h52 : rvCrc[28] <= 32'hbc924678;
8'h53 : rvCrc[28] <= 32'hc92c00cf;
8'h54 : rvCrc[28] <= 32'h85d6cc7d;
8'h55 : rvCrc[28] <= 32'hf0688aca;
8'h56 : rvCrc[28] <= 32'h6eaa4113;
8'h57 : rvCrc[28] <= 32'h1b1407a4;
8'h58 : rvCrc[28] <= 32'hf75fd877;
8'h59 : rvCrc[28] <= 32'h82e19ec0;
8'h5a : rvCrc[28] <= 32'h1c235519;
8'h5b : rvCrc[28] <= 32'h699d13ae;
8'h5c : rvCrc[28] <= 32'h2567df1c;
8'h5d : rvCrc[28] <= 32'h50d999ab;
8'h5e : rvCrc[28] <= 32'hce1b5272;
8'h5f : rvCrc[28] <= 32'hbba514c5;
8'h60 : rvCrc[28] <= 32'h990b8689;
8'h61 : rvCrc[28] <= 32'hecb5c03e;
8'h62 : rvCrc[28] <= 32'h72770be7;
8'h63 : rvCrc[28] <= 32'h07c94d50;
8'h64 : rvCrc[28] <= 32'h4b3381e2;
8'h65 : rvCrc[28] <= 32'h3e8dc755;
8'h66 : rvCrc[28] <= 32'ha04f0c8c;
8'h67 : rvCrc[28] <= 32'hd5f14a3b;
8'h68 : rvCrc[28] <= 32'h39ba95e8;
8'h69 : rvCrc[28] <= 32'h4c04d35f;
8'h6a : rvCrc[28] <= 32'hd2c61886;
8'h6b : rvCrc[28] <= 32'ha7785e31;
8'h6c : rvCrc[28] <= 32'heb829283;
8'h6d : rvCrc[28] <= 32'h9e3cd434;
8'h6e : rvCrc[28] <= 32'h00fe1fed;
8'h6f : rvCrc[28] <= 32'h7540595a;
8'h70 : rvCrc[28] <= 32'hdca8bdfc;
8'h71 : rvCrc[28] <= 32'ha916fb4b;
8'h72 : rvCrc[28] <= 32'h37d43092;
8'h73 : rvCrc[28] <= 32'h426a7625;
8'h74 : rvCrc[28] <= 32'h0e90ba97;
8'h75 : rvCrc[28] <= 32'h7b2efc20;
8'h76 : rvCrc[28] <= 32'he5ec37f9;
8'h77 : rvCrc[28] <= 32'h9052714e;
8'h78 : rvCrc[28] <= 32'h7c19ae9d;
8'h79 : rvCrc[28] <= 32'h09a7e82a;
8'h7a : rvCrc[28] <= 32'h976523f3;
8'h7b : rvCrc[28] <= 32'he2db6544;
8'h7c : rvCrc[28] <= 32'hae21a9f6;
8'h7d : rvCrc[28] <= 32'hdb9fef41;
8'h7e : rvCrc[28] <= 32'h455d2498;
8'h7f : rvCrc[28] <= 32'h30e3622f;
8'h80 : rvCrc[28] <= 32'h249be0c6;
8'h81 : rvCrc[28] <= 32'h5125a671;
8'h82 : rvCrc[28] <= 32'hcfe76da8;
8'h83 : rvCrc[28] <= 32'hba592b1f;
8'h84 : rvCrc[28] <= 32'hf6a3e7ad;
8'h85 : rvCrc[28] <= 32'h831da11a;
8'h86 : rvCrc[28] <= 32'h1ddf6ac3;
8'h87 : rvCrc[28] <= 32'h68612c74;
8'h88 : rvCrc[28] <= 32'h842af3a7;
8'h89 : rvCrc[28] <= 32'hf194b510;
8'h8a : rvCrc[28] <= 32'h6f567ec9;
8'h8b : rvCrc[28] <= 32'h1ae8387e;
8'h8c : rvCrc[28] <= 32'h5612f4cc;
8'h8d : rvCrc[28] <= 32'h23acb27b;
8'h8e : rvCrc[28] <= 32'hbd6e79a2;
8'h8f : rvCrc[28] <= 32'hc8d03f15;
8'h90 : rvCrc[28] <= 32'h6138dbb3;
8'h91 : rvCrc[28] <= 32'h14869d04;
8'h92 : rvCrc[28] <= 32'h8a4456dd;
8'h93 : rvCrc[28] <= 32'hfffa106a;
8'h94 : rvCrc[28] <= 32'hb300dcd8;
8'h95 : rvCrc[28] <= 32'hc6be9a6f;
8'h96 : rvCrc[28] <= 32'h587c51b6;
8'h97 : rvCrc[28] <= 32'h2dc21701;
8'h98 : rvCrc[28] <= 32'hc189c8d2;
8'h99 : rvCrc[28] <= 32'hb4378e65;
8'h9a : rvCrc[28] <= 32'h2af545bc;
8'h9b : rvCrc[28] <= 32'h5f4b030b;
8'h9c : rvCrc[28] <= 32'h13b1cfb9;
8'h9d : rvCrc[28] <= 32'h660f890e;
8'h9e : rvCrc[28] <= 32'hf8cd42d7;
8'h9f : rvCrc[28] <= 32'h8d730460;
8'ha0 : rvCrc[28] <= 32'hafdd962c;
8'ha1 : rvCrc[28] <= 32'hda63d09b;
8'ha2 : rvCrc[28] <= 32'h44a11b42;
8'ha3 : rvCrc[28] <= 32'h311f5df5;
8'ha4 : rvCrc[28] <= 32'h7de59147;
8'ha5 : rvCrc[28] <= 32'h085bd7f0;
8'ha6 : rvCrc[28] <= 32'h96991c29;
8'ha7 : rvCrc[28] <= 32'he3275a9e;
8'ha8 : rvCrc[28] <= 32'h0f6c854d;
8'ha9 : rvCrc[28] <= 32'h7ad2c3fa;
8'haa : rvCrc[28] <= 32'he4100823;
8'hab : rvCrc[28] <= 32'h91ae4e94;
8'hac : rvCrc[28] <= 32'hdd548226;
8'had : rvCrc[28] <= 32'ha8eac491;
8'hae : rvCrc[28] <= 32'h36280f48;
8'haf : rvCrc[28] <= 32'h439649ff;
8'hb0 : rvCrc[28] <= 32'hea7ead59;
8'hb1 : rvCrc[28] <= 32'h9fc0ebee;
8'hb2 : rvCrc[28] <= 32'h01022037;
8'hb3 : rvCrc[28] <= 32'h74bc6680;
8'hb4 : rvCrc[28] <= 32'h3846aa32;
8'hb5 : rvCrc[28] <= 32'h4df8ec85;
8'hb6 : rvCrc[28] <= 32'hd33a275c;
8'hb7 : rvCrc[28] <= 32'ha68461eb;
8'hb8 : rvCrc[28] <= 32'h4acfbe38;
8'hb9 : rvCrc[28] <= 32'h3f71f88f;
8'hba : rvCrc[28] <= 32'ha1b33356;
8'hbb : rvCrc[28] <= 32'hd40d75e1;
8'hbc : rvCrc[28] <= 32'h98f7b953;
8'hbd : rvCrc[28] <= 32'hed49ffe4;
8'hbe : rvCrc[28] <= 32'h738b343d;
8'hbf : rvCrc[28] <= 32'h0635728a;
8'hc0 : rvCrc[28] <= 32'h36d610a5;
8'hc1 : rvCrc[28] <= 32'h43685612;
8'hc2 : rvCrc[28] <= 32'hddaa9dcb;
8'hc3 : rvCrc[28] <= 32'ha814db7c;
8'hc4 : rvCrc[28] <= 32'he4ee17ce;
8'hc5 : rvCrc[28] <= 32'h91505179;
8'hc6 : rvCrc[28] <= 32'h0f929aa0;
8'hc7 : rvCrc[28] <= 32'h7a2cdc17;
8'hc8 : rvCrc[28] <= 32'h966703c4;
8'hc9 : rvCrc[28] <= 32'he3d94573;
8'hca : rvCrc[28] <= 32'h7d1b8eaa;
8'hcb : rvCrc[28] <= 32'h08a5c81d;
8'hcc : rvCrc[28] <= 32'h445f04af;
8'hcd : rvCrc[28] <= 32'h31e14218;
8'hce : rvCrc[28] <= 32'haf2389c1;
8'hcf : rvCrc[28] <= 32'hda9dcf76;
8'hd0 : rvCrc[28] <= 32'h73752bd0;
8'hd1 : rvCrc[28] <= 32'h06cb6d67;
8'hd2 : rvCrc[28] <= 32'h9809a6be;
8'hd3 : rvCrc[28] <= 32'hedb7e009;
8'hd4 : rvCrc[28] <= 32'ha14d2cbb;
8'hd5 : rvCrc[28] <= 32'hd4f36a0c;
8'hd6 : rvCrc[28] <= 32'h4a31a1d5;
8'hd7 : rvCrc[28] <= 32'h3f8fe762;
8'hd8 : rvCrc[28] <= 32'hd3c438b1;
8'hd9 : rvCrc[28] <= 32'ha67a7e06;
8'hda : rvCrc[28] <= 32'h38b8b5df;
8'hdb : rvCrc[28] <= 32'h4d06f368;
8'hdc : rvCrc[28] <= 32'h01fc3fda;
8'hdd : rvCrc[28] <= 32'h7442796d;
8'hde : rvCrc[28] <= 32'hea80b2b4;
8'hdf : rvCrc[28] <= 32'h9f3ef403;
8'he0 : rvCrc[28] <= 32'hbd90664f;
8'he1 : rvCrc[28] <= 32'hc82e20f8;
8'he2 : rvCrc[28] <= 32'h56eceb21;
8'he3 : rvCrc[28] <= 32'h2352ad96;
8'he4 : rvCrc[28] <= 32'h6fa86124;
8'he5 : rvCrc[28] <= 32'h1a162793;
8'he6 : rvCrc[28] <= 32'h84d4ec4a;
8'he7 : rvCrc[28] <= 32'hf16aaafd;
8'he8 : rvCrc[28] <= 32'h1d21752e;
8'he9 : rvCrc[28] <= 32'h689f3399;
8'hea : rvCrc[28] <= 32'hf65df840;
8'heb : rvCrc[28] <= 32'h83e3bef7;
8'hec : rvCrc[28] <= 32'hcf197245;
8'hed : rvCrc[28] <= 32'hbaa734f2;
8'hee : rvCrc[28] <= 32'h2465ff2b;
8'hef : rvCrc[28] <= 32'h51dbb99c;
8'hf0 : rvCrc[28] <= 32'hf8335d3a;
8'hf1 : rvCrc[28] <= 32'h8d8d1b8d;
8'hf2 : rvCrc[28] <= 32'h134fd054;
8'hf3 : rvCrc[28] <= 32'h66f196e3;
8'hf4 : rvCrc[28] <= 32'h2a0b5a51;
8'hf5 : rvCrc[28] <= 32'h5fb51ce6;
8'hf6 : rvCrc[28] <= 32'hc177d73f;
8'hf7 : rvCrc[28] <= 32'hb4c99188;
8'hf8 : rvCrc[28] <= 32'h58824e5b;
8'hf9 : rvCrc[28] <= 32'h2d3c08ec;
8'hfa : rvCrc[28] <= 32'hb3fec335;
8'hfb : rvCrc[28] <= 32'hc6408582;
8'hfc : rvCrc[28] <= 32'h8aba4930;
8'hfd : rvCrc[28] <= 32'hff040f87;
8'hfe : rvCrc[28] <= 32'h61c6c45e;
8'hff : rvCrc[28] <= 32'h147882e9;
endcase
case(iv_Input[239:232])
8'h00 : rvCrc[29] <= 32'h00000000;
8'h01 : rvCrc[29] <= 32'h4937c18c;
8'h02 : rvCrc[29] <= 32'h926f8318;
8'h03 : rvCrc[29] <= 32'hdb584294;
8'h04 : rvCrc[29] <= 32'h201e1b87;
8'h05 : rvCrc[29] <= 32'h6929da0b;
8'h06 : rvCrc[29] <= 32'hb271989f;
8'h07 : rvCrc[29] <= 32'hfb465913;
8'h08 : rvCrc[29] <= 32'h403c370e;
8'h09 : rvCrc[29] <= 32'h090bf682;
8'h0a : rvCrc[29] <= 32'hd253b416;
8'h0b : rvCrc[29] <= 32'h9b64759a;
8'h0c : rvCrc[29] <= 32'h60222c89;
8'h0d : rvCrc[29] <= 32'h2915ed05;
8'h0e : rvCrc[29] <= 32'hf24daf91;
8'h0f : rvCrc[29] <= 32'hbb7a6e1d;
8'h10 : rvCrc[29] <= 32'h80786e1c;
8'h11 : rvCrc[29] <= 32'hc94faf90;
8'h12 : rvCrc[29] <= 32'h1217ed04;
8'h13 : rvCrc[29] <= 32'h5b202c88;
8'h14 : rvCrc[29] <= 32'ha066759b;
8'h15 : rvCrc[29] <= 32'he951b417;
8'h16 : rvCrc[29] <= 32'h3209f683;
8'h17 : rvCrc[29] <= 32'h7b3e370f;
8'h18 : rvCrc[29] <= 32'hc0445912;
8'h19 : rvCrc[29] <= 32'h8973989e;
8'h1a : rvCrc[29] <= 32'h522bda0a;
8'h1b : rvCrc[29] <= 32'h1b1c1b86;
8'h1c : rvCrc[29] <= 32'he05a4295;
8'h1d : rvCrc[29] <= 32'ha96d8319;
8'h1e : rvCrc[29] <= 32'h7235c18d;
8'h1f : rvCrc[29] <= 32'h3b020001;
8'h20 : rvCrc[29] <= 32'h0431c18f;
8'h21 : rvCrc[29] <= 32'h4d060003;
8'h22 : rvCrc[29] <= 32'h965e4297;
8'h23 : rvCrc[29] <= 32'hdf69831b;
8'h24 : rvCrc[29] <= 32'h242fda08;
8'h25 : rvCrc[29] <= 32'h6d181b84;
8'h26 : rvCrc[29] <= 32'hb6405910;
8'h27 : rvCrc[29] <= 32'hff77989c;
8'h28 : rvCrc[29] <= 32'h440df681;
8'h29 : rvCrc[29] <= 32'h0d3a370d;
8'h2a : rvCrc[29] <= 32'hd6627599;
8'h2b : rvCrc[29] <= 32'h9f55b415;
8'h2c : rvCrc[29] <= 32'h6413ed06;
8'h2d : rvCrc[29] <= 32'h2d242c8a;
8'h2e : rvCrc[29] <= 32'hf67c6e1e;
8'h2f : rvCrc[29] <= 32'hbf4baf92;
8'h30 : rvCrc[29] <= 32'h8449af93;
8'h31 : rvCrc[29] <= 32'hcd7e6e1f;
8'h32 : rvCrc[29] <= 32'h16262c8b;
8'h33 : rvCrc[29] <= 32'h5f11ed07;
8'h34 : rvCrc[29] <= 32'ha457b414;
8'h35 : rvCrc[29] <= 32'hed607598;
8'h36 : rvCrc[29] <= 32'h3638370c;
8'h37 : rvCrc[29] <= 32'h7f0ff680;
8'h38 : rvCrc[29] <= 32'hc475989d;
8'h39 : rvCrc[29] <= 32'h8d425911;
8'h3a : rvCrc[29] <= 32'h561a1b85;
8'h3b : rvCrc[29] <= 32'h1f2dda09;
8'h3c : rvCrc[29] <= 32'he46b831a;
8'h3d : rvCrc[29] <= 32'had5c4296;
8'h3e : rvCrc[29] <= 32'h76040002;
8'h3f : rvCrc[29] <= 32'h3f33c18e;
8'h40 : rvCrc[29] <= 32'h0863831e;
8'h41 : rvCrc[29] <= 32'h41544292;
8'h42 : rvCrc[29] <= 32'h9a0c0006;
8'h43 : rvCrc[29] <= 32'hd33bc18a;
8'h44 : rvCrc[29] <= 32'h287d9899;
8'h45 : rvCrc[29] <= 32'h614a5915;
8'h46 : rvCrc[29] <= 32'hba121b81;
8'h47 : rvCrc[29] <= 32'hf325da0d;
8'h48 : rvCrc[29] <= 32'h485fb410;
8'h49 : rvCrc[29] <= 32'h0168759c;
8'h4a : rvCrc[29] <= 32'hda303708;
8'h4b : rvCrc[29] <= 32'h9307f684;
8'h4c : rvCrc[29] <= 32'h6841af97;
8'h4d : rvCrc[29] <= 32'h21766e1b;
8'h4e : rvCrc[29] <= 32'hfa2e2c8f;
8'h4f : rvCrc[29] <= 32'hb319ed03;
8'h50 : rvCrc[29] <= 32'h881bed02;
8'h51 : rvCrc[29] <= 32'hc12c2c8e;
8'h52 : rvCrc[29] <= 32'h1a746e1a;
8'h53 : rvCrc[29] <= 32'h5343af96;
8'h54 : rvCrc[29] <= 32'ha805f685;
8'h55 : rvCrc[29] <= 32'he1323709;
8'h56 : rvCrc[29] <= 32'h3a6a759d;
8'h57 : rvCrc[29] <= 32'h735db411;
8'h58 : rvCrc[29] <= 32'hc827da0c;
8'h59 : rvCrc[29] <= 32'h81101b80;
8'h5a : rvCrc[29] <= 32'h5a485914;
8'h5b : rvCrc[29] <= 32'h137f9898;
8'h5c : rvCrc[29] <= 32'he839c18b;
8'h5d : rvCrc[29] <= 32'ha10e0007;
8'h5e : rvCrc[29] <= 32'h7a564293;
8'h5f : rvCrc[29] <= 32'h3361831f;
8'h60 : rvCrc[29] <= 32'h0c524291;
8'h61 : rvCrc[29] <= 32'h4565831d;
8'h62 : rvCrc[29] <= 32'h9e3dc189;
8'h63 : rvCrc[29] <= 32'hd70a0005;
8'h64 : rvCrc[29] <= 32'h2c4c5916;
8'h65 : rvCrc[29] <= 32'h657b989a;
8'h66 : rvCrc[29] <= 32'hbe23da0e;
8'h67 : rvCrc[29] <= 32'hf7141b82;
8'h68 : rvCrc[29] <= 32'h4c6e759f;
8'h69 : rvCrc[29] <= 32'h0559b413;
8'h6a : rvCrc[29] <= 32'hde01f687;
8'h6b : rvCrc[29] <= 32'h9736370b;
8'h6c : rvCrc[29] <= 32'h6c706e18;
8'h6d : rvCrc[29] <= 32'h2547af94;
8'h6e : rvCrc[29] <= 32'hfe1fed00;
8'h6f : rvCrc[29] <= 32'hb7282c8c;
8'h70 : rvCrc[29] <= 32'h8c2a2c8d;
8'h71 : rvCrc[29] <= 32'hc51ded01;
8'h72 : rvCrc[29] <= 32'h1e45af95;
8'h73 : rvCrc[29] <= 32'h57726e19;
8'h74 : rvCrc[29] <= 32'hac34370a;
8'h75 : rvCrc[29] <= 32'he503f686;
8'h76 : rvCrc[29] <= 32'h3e5bb412;
8'h77 : rvCrc[29] <= 32'h776c759e;
8'h78 : rvCrc[29] <= 32'hcc161b83;
8'h79 : rvCrc[29] <= 32'h8521da0f;
8'h7a : rvCrc[29] <= 32'h5e79989b;
8'h7b : rvCrc[29] <= 32'h174e5917;
8'h7c : rvCrc[29] <= 32'hec080004;
8'h7d : rvCrc[29] <= 32'ha53fc188;
8'h7e : rvCrc[29] <= 32'h7e67831c;
8'h7f : rvCrc[29] <= 32'h37504290;
8'h80 : rvCrc[29] <= 32'h10c7063c;
8'h81 : rvCrc[29] <= 32'h59f0c7b0;
8'h82 : rvCrc[29] <= 32'h82a88524;
8'h83 : rvCrc[29] <= 32'hcb9f44a8;
8'h84 : rvCrc[29] <= 32'h30d91dbb;
8'h85 : rvCrc[29] <= 32'h79eedc37;
8'h86 : rvCrc[29] <= 32'ha2b69ea3;
8'h87 : rvCrc[29] <= 32'heb815f2f;
8'h88 : rvCrc[29] <= 32'h50fb3132;
8'h89 : rvCrc[29] <= 32'h19ccf0be;
8'h8a : rvCrc[29] <= 32'hc294b22a;
8'h8b : rvCrc[29] <= 32'h8ba373a6;
8'h8c : rvCrc[29] <= 32'h70e52ab5;
8'h8d : rvCrc[29] <= 32'h39d2eb39;
8'h8e : rvCrc[29] <= 32'he28aa9ad;
8'h8f : rvCrc[29] <= 32'habbd6821;
8'h90 : rvCrc[29] <= 32'h90bf6820;
8'h91 : rvCrc[29] <= 32'hd988a9ac;
8'h92 : rvCrc[29] <= 32'h02d0eb38;
8'h93 : rvCrc[29] <= 32'h4be72ab4;
8'h94 : rvCrc[29] <= 32'hb0a173a7;
8'h95 : rvCrc[29] <= 32'hf996b22b;
8'h96 : rvCrc[29] <= 32'h22cef0bf;
8'h97 : rvCrc[29] <= 32'h6bf93133;
8'h98 : rvCrc[29] <= 32'hd0835f2e;
8'h99 : rvCrc[29] <= 32'h99b49ea2;
8'h9a : rvCrc[29] <= 32'h42ecdc36;
8'h9b : rvCrc[29] <= 32'h0bdb1dba;
8'h9c : rvCrc[29] <= 32'hf09d44a9;
8'h9d : rvCrc[29] <= 32'hb9aa8525;
8'h9e : rvCrc[29] <= 32'h62f2c7b1;
8'h9f : rvCrc[29] <= 32'h2bc5063d;
8'ha0 : rvCrc[29] <= 32'h14f6c7b3;
8'ha1 : rvCrc[29] <= 32'h5dc1063f;
8'ha2 : rvCrc[29] <= 32'h869944ab;
8'ha3 : rvCrc[29] <= 32'hcfae8527;
8'ha4 : rvCrc[29] <= 32'h34e8dc34;
8'ha5 : rvCrc[29] <= 32'h7ddf1db8;
8'ha6 : rvCrc[29] <= 32'ha6875f2c;
8'ha7 : rvCrc[29] <= 32'hefb09ea0;
8'ha8 : rvCrc[29] <= 32'h54caf0bd;
8'ha9 : rvCrc[29] <= 32'h1dfd3131;
8'haa : rvCrc[29] <= 32'hc6a573a5;
8'hab : rvCrc[29] <= 32'h8f92b229;
8'hac : rvCrc[29] <= 32'h74d4eb3a;
8'had : rvCrc[29] <= 32'h3de32ab6;
8'hae : rvCrc[29] <= 32'he6bb6822;
8'haf : rvCrc[29] <= 32'haf8ca9ae;
8'hb0 : rvCrc[29] <= 32'h948ea9af;
8'hb1 : rvCrc[29] <= 32'hddb96823;
8'hb2 : rvCrc[29] <= 32'h06e12ab7;
8'hb3 : rvCrc[29] <= 32'h4fd6eb3b;
8'hb4 : rvCrc[29] <= 32'hb490b228;
8'hb5 : rvCrc[29] <= 32'hfda773a4;
8'hb6 : rvCrc[29] <= 32'h26ff3130;
8'hb7 : rvCrc[29] <= 32'h6fc8f0bc;
8'hb8 : rvCrc[29] <= 32'hd4b29ea1;
8'hb9 : rvCrc[29] <= 32'h9d855f2d;
8'hba : rvCrc[29] <= 32'h46dd1db9;
8'hbb : rvCrc[29] <= 32'h0feadc35;
8'hbc : rvCrc[29] <= 32'hf4ac8526;
8'hbd : rvCrc[29] <= 32'hbd9b44aa;
8'hbe : rvCrc[29] <= 32'h66c3063e;
8'hbf : rvCrc[29] <= 32'h2ff4c7b2;
8'hc0 : rvCrc[29] <= 32'h18a48522;
8'hc1 : rvCrc[29] <= 32'h519344ae;
8'hc2 : rvCrc[29] <= 32'h8acb063a;
8'hc3 : rvCrc[29] <= 32'hc3fcc7b6;
8'hc4 : rvCrc[29] <= 32'h38ba9ea5;
8'hc5 : rvCrc[29] <= 32'h718d5f29;
8'hc6 : rvCrc[29] <= 32'haad51dbd;
8'hc7 : rvCrc[29] <= 32'he3e2dc31;
8'hc8 : rvCrc[29] <= 32'h5898b22c;
8'hc9 : rvCrc[29] <= 32'h11af73a0;
8'hca : rvCrc[29] <= 32'hcaf73134;
8'hcb : rvCrc[29] <= 32'h83c0f0b8;
8'hcc : rvCrc[29] <= 32'h7886a9ab;
8'hcd : rvCrc[29] <= 32'h31b16827;
8'hce : rvCrc[29] <= 32'heae92ab3;
8'hcf : rvCrc[29] <= 32'ha3deeb3f;
8'hd0 : rvCrc[29] <= 32'h98dceb3e;
8'hd1 : rvCrc[29] <= 32'hd1eb2ab2;
8'hd2 : rvCrc[29] <= 32'h0ab36826;
8'hd3 : rvCrc[29] <= 32'h4384a9aa;
8'hd4 : rvCrc[29] <= 32'hb8c2f0b9;
8'hd5 : rvCrc[29] <= 32'hf1f53135;
8'hd6 : rvCrc[29] <= 32'h2aad73a1;
8'hd7 : rvCrc[29] <= 32'h639ab22d;
8'hd8 : rvCrc[29] <= 32'hd8e0dc30;
8'hd9 : rvCrc[29] <= 32'h91d71dbc;
8'hda : rvCrc[29] <= 32'h4a8f5f28;
8'hdb : rvCrc[29] <= 32'h03b89ea4;
8'hdc : rvCrc[29] <= 32'hf8fec7b7;
8'hdd : rvCrc[29] <= 32'hb1c9063b;
8'hde : rvCrc[29] <= 32'h6a9144af;
8'hdf : rvCrc[29] <= 32'h23a68523;
8'he0 : rvCrc[29] <= 32'h1c9544ad;
8'he1 : rvCrc[29] <= 32'h55a28521;
8'he2 : rvCrc[29] <= 32'h8efac7b5;
8'he3 : rvCrc[29] <= 32'hc7cd0639;
8'he4 : rvCrc[29] <= 32'h3c8b5f2a;
8'he5 : rvCrc[29] <= 32'h75bc9ea6;
8'he6 : rvCrc[29] <= 32'haee4dc32;
8'he7 : rvCrc[29] <= 32'he7d31dbe;
8'he8 : rvCrc[29] <= 32'h5ca973a3;
8'he9 : rvCrc[29] <= 32'h159eb22f;
8'hea : rvCrc[29] <= 32'hcec6f0bb;
8'heb : rvCrc[29] <= 32'h87f13137;
8'hec : rvCrc[29] <= 32'h7cb76824;
8'hed : rvCrc[29] <= 32'h3580a9a8;
8'hee : rvCrc[29] <= 32'heed8eb3c;
8'hef : rvCrc[29] <= 32'ha7ef2ab0;
8'hf0 : rvCrc[29] <= 32'h9ced2ab1;
8'hf1 : rvCrc[29] <= 32'hd5daeb3d;
8'hf2 : rvCrc[29] <= 32'h0e82a9a9;
8'hf3 : rvCrc[29] <= 32'h47b56825;
8'hf4 : rvCrc[29] <= 32'hbcf33136;
8'hf5 : rvCrc[29] <= 32'hf5c4f0ba;
8'hf6 : rvCrc[29] <= 32'h2e9cb22e;
8'hf7 : rvCrc[29] <= 32'h67ab73a2;
8'hf8 : rvCrc[29] <= 32'hdcd11dbf;
8'hf9 : rvCrc[29] <= 32'h95e6dc33;
8'hfa : rvCrc[29] <= 32'h4ebe9ea7;
8'hfb : rvCrc[29] <= 32'h07895f2b;
8'hfc : rvCrc[29] <= 32'hfccf0638;
8'hfd : rvCrc[29] <= 32'hb5f8c7b4;
8'hfe : rvCrc[29] <= 32'h6ea08520;
8'hff : rvCrc[29] <= 32'h279744ac;
endcase
case(iv_Input[247:240])
8'h00 : rvCrc[30] <= 32'h00000000;
8'h01 : rvCrc[30] <= 32'h218e0c78;
8'h02 : rvCrc[30] <= 32'h431c18f0;
8'h03 : rvCrc[30] <= 32'h62921488;
8'h04 : rvCrc[30] <= 32'h863831e0;
8'h05 : rvCrc[30] <= 32'ha7b63d98;
8'h06 : rvCrc[30] <= 32'hc5242910;
8'h07 : rvCrc[30] <= 32'he4aa2568;
8'h08 : rvCrc[30] <= 32'h08b17e77;
8'h09 : rvCrc[30] <= 32'h293f720f;
8'h0a : rvCrc[30] <= 32'h4bad6687;
8'h0b : rvCrc[30] <= 32'h6a236aff;
8'h0c : rvCrc[30] <= 32'h8e894f97;
8'h0d : rvCrc[30] <= 32'haf0743ef;
8'h0e : rvCrc[30] <= 32'hcd955767;
8'h0f : rvCrc[30] <= 32'hec1b5b1f;
8'h10 : rvCrc[30] <= 32'h1162fcee;
8'h11 : rvCrc[30] <= 32'h30ecf096;
8'h12 : rvCrc[30] <= 32'h527ee41e;
8'h13 : rvCrc[30] <= 32'h73f0e866;
8'h14 : rvCrc[30] <= 32'h975acd0e;
8'h15 : rvCrc[30] <= 32'hb6d4c176;
8'h16 : rvCrc[30] <= 32'hd446d5fe;
8'h17 : rvCrc[30] <= 32'hf5c8d986;
8'h18 : rvCrc[30] <= 32'h19d38299;
8'h19 : rvCrc[30] <= 32'h385d8ee1;
8'h1a : rvCrc[30] <= 32'h5acf9a69;
8'h1b : rvCrc[30] <= 32'h7b419611;
8'h1c : rvCrc[30] <= 32'h9febb379;
8'h1d : rvCrc[30] <= 32'hbe65bf01;
8'h1e : rvCrc[30] <= 32'hdcf7ab89;
8'h1f : rvCrc[30] <= 32'hfd79a7f1;
8'h20 : rvCrc[30] <= 32'h22c5f9dc;
8'h21 : rvCrc[30] <= 32'h034bf5a4;
8'h22 : rvCrc[30] <= 32'h61d9e12c;
8'h23 : rvCrc[30] <= 32'h4057ed54;
8'h24 : rvCrc[30] <= 32'ha4fdc83c;
8'h25 : rvCrc[30] <= 32'h8573c444;
8'h26 : rvCrc[30] <= 32'he7e1d0cc;
8'h27 : rvCrc[30] <= 32'hc66fdcb4;
8'h28 : rvCrc[30] <= 32'h2a7487ab;
8'h29 : rvCrc[30] <= 32'h0bfa8bd3;
8'h2a : rvCrc[30] <= 32'h69689f5b;
8'h2b : rvCrc[30] <= 32'h48e69323;
8'h2c : rvCrc[30] <= 32'hac4cb64b;
8'h2d : rvCrc[30] <= 32'h8dc2ba33;
8'h2e : rvCrc[30] <= 32'hef50aebb;
8'h2f : rvCrc[30] <= 32'hcedea2c3;
8'h30 : rvCrc[30] <= 32'h33a70532;
8'h31 : rvCrc[30] <= 32'h1229094a;
8'h32 : rvCrc[30] <= 32'h70bb1dc2;
8'h33 : rvCrc[30] <= 32'h513511ba;
8'h34 : rvCrc[30] <= 32'hb59f34d2;
8'h35 : rvCrc[30] <= 32'h941138aa;
8'h36 : rvCrc[30] <= 32'hf6832c22;
8'h37 : rvCrc[30] <= 32'hd70d205a;
8'h38 : rvCrc[30] <= 32'h3b167b45;
8'h39 : rvCrc[30] <= 32'h1a98773d;
8'h3a : rvCrc[30] <= 32'h780a63b5;
8'h3b : rvCrc[30] <= 32'h59846fcd;
8'h3c : rvCrc[30] <= 32'hbd2e4aa5;
8'h3d : rvCrc[30] <= 32'h9ca046dd;
8'h3e : rvCrc[30] <= 32'hfe325255;
8'h3f : rvCrc[30] <= 32'hdfbc5e2d;
8'h40 : rvCrc[30] <= 32'h458bf3b8;
8'h41 : rvCrc[30] <= 32'h6405ffc0;
8'h42 : rvCrc[30] <= 32'h0697eb48;
8'h43 : rvCrc[30] <= 32'h2719e730;
8'h44 : rvCrc[30] <= 32'hc3b3c258;
8'h45 : rvCrc[30] <= 32'he23dce20;
8'h46 : rvCrc[30] <= 32'h80afdaa8;
8'h47 : rvCrc[30] <= 32'ha121d6d0;
8'h48 : rvCrc[30] <= 32'h4d3a8dcf;
8'h49 : rvCrc[30] <= 32'h6cb481b7;
8'h4a : rvCrc[30] <= 32'h0e26953f;
8'h4b : rvCrc[30] <= 32'h2fa89947;
8'h4c : rvCrc[30] <= 32'hcb02bc2f;
8'h4d : rvCrc[30] <= 32'hea8cb057;
8'h4e : rvCrc[30] <= 32'h881ea4df;
8'h4f : rvCrc[30] <= 32'ha990a8a7;
8'h50 : rvCrc[30] <= 32'h54e90f56;
8'h51 : rvCrc[30] <= 32'h7567032e;
8'h52 : rvCrc[30] <= 32'h17f517a6;
8'h53 : rvCrc[30] <= 32'h367b1bde;
8'h54 : rvCrc[30] <= 32'hd2d13eb6;
8'h55 : rvCrc[30] <= 32'hf35f32ce;
8'h56 : rvCrc[30] <= 32'h91cd2646;
8'h57 : rvCrc[30] <= 32'hb0432a3e;
8'h58 : rvCrc[30] <= 32'h5c587121;
8'h59 : rvCrc[30] <= 32'h7dd67d59;
8'h5a : rvCrc[30] <= 32'h1f4469d1;
8'h5b : rvCrc[30] <= 32'h3eca65a9;
8'h5c : rvCrc[30] <= 32'hda6040c1;
8'h5d : rvCrc[30] <= 32'hfbee4cb9;
8'h5e : rvCrc[30] <= 32'h997c5831;
8'h5f : rvCrc[30] <= 32'hb8f25449;
8'h60 : rvCrc[30] <= 32'h674e0a64;
8'h61 : rvCrc[30] <= 32'h46c0061c;
8'h62 : rvCrc[30] <= 32'h24521294;
8'h63 : rvCrc[30] <= 32'h05dc1eec;
8'h64 : rvCrc[30] <= 32'he1763b84;
8'h65 : rvCrc[30] <= 32'hc0f837fc;
8'h66 : rvCrc[30] <= 32'ha26a2374;
8'h67 : rvCrc[30] <= 32'h83e42f0c;
8'h68 : rvCrc[30] <= 32'h6fff7413;
8'h69 : rvCrc[30] <= 32'h4e71786b;
8'h6a : rvCrc[30] <= 32'h2ce36ce3;
8'h6b : rvCrc[30] <= 32'h0d6d609b;
8'h6c : rvCrc[30] <= 32'he9c745f3;
8'h6d : rvCrc[30] <= 32'hc849498b;
8'h6e : rvCrc[30] <= 32'haadb5d03;
8'h6f : rvCrc[30] <= 32'h8b55517b;
8'h70 : rvCrc[30] <= 32'h762cf68a;
8'h71 : rvCrc[30] <= 32'h57a2faf2;
8'h72 : rvCrc[30] <= 32'h3530ee7a;
8'h73 : rvCrc[30] <= 32'h14bee202;
8'h74 : rvCrc[30] <= 32'hf014c76a;
8'h75 : rvCrc[30] <= 32'hd19acb12;
8'h76 : rvCrc[30] <= 32'hb308df9a;
8'h77 : rvCrc[30] <= 32'h9286d3e2;
8'h78 : rvCrc[30] <= 32'h7e9d88fd;
8'h79 : rvCrc[30] <= 32'h5f138485;
8'h7a : rvCrc[30] <= 32'h3d81900d;
8'h7b : rvCrc[30] <= 32'h1c0f9c75;
8'h7c : rvCrc[30] <= 32'hf8a5b91d;
8'h7d : rvCrc[30] <= 32'hd92bb565;
8'h7e : rvCrc[30] <= 32'hbbb9a1ed;
8'h7f : rvCrc[30] <= 32'h9a37ad95;
8'h80 : rvCrc[30] <= 32'h8b17e770;
8'h81 : rvCrc[30] <= 32'haa99eb08;
8'h82 : rvCrc[30] <= 32'hc80bff80;
8'h83 : rvCrc[30] <= 32'he985f3f8;
8'h84 : rvCrc[30] <= 32'h0d2fd690;
8'h85 : rvCrc[30] <= 32'h2ca1dae8;
8'h86 : rvCrc[30] <= 32'h4e33ce60;
8'h87 : rvCrc[30] <= 32'h6fbdc218;
8'h88 : rvCrc[30] <= 32'h83a69907;
8'h89 : rvCrc[30] <= 32'ha228957f;
8'h8a : rvCrc[30] <= 32'hc0ba81f7;
8'h8b : rvCrc[30] <= 32'he1348d8f;
8'h8c : rvCrc[30] <= 32'h059ea8e7;
8'h8d : rvCrc[30] <= 32'h2410a49f;
8'h8e : rvCrc[30] <= 32'h4682b017;
8'h8f : rvCrc[30] <= 32'h670cbc6f;
8'h90 : rvCrc[30] <= 32'h9a751b9e;
8'h91 : rvCrc[30] <= 32'hbbfb17e6;
8'h92 : rvCrc[30] <= 32'hd969036e;
8'h93 : rvCrc[30] <= 32'hf8e70f16;
8'h94 : rvCrc[30] <= 32'h1c4d2a7e;
8'h95 : rvCrc[30] <= 32'h3dc32606;
8'h96 : rvCrc[30] <= 32'h5f51328e;
8'h97 : rvCrc[30] <= 32'h7edf3ef6;
8'h98 : rvCrc[30] <= 32'h92c465e9;
8'h99 : rvCrc[30] <= 32'hb34a6991;
8'h9a : rvCrc[30] <= 32'hd1d87d19;
8'h9b : rvCrc[30] <= 32'hf0567161;
8'h9c : rvCrc[30] <= 32'h14fc5409;
8'h9d : rvCrc[30] <= 32'h35725871;
8'h9e : rvCrc[30] <= 32'h57e04cf9;
8'h9f : rvCrc[30] <= 32'h766e4081;
8'ha0 : rvCrc[30] <= 32'ha9d21eac;
8'ha1 : rvCrc[30] <= 32'h885c12d4;
8'ha2 : rvCrc[30] <= 32'heace065c;
8'ha3 : rvCrc[30] <= 32'hcb400a24;
8'ha4 : rvCrc[30] <= 32'h2fea2f4c;
8'ha5 : rvCrc[30] <= 32'h0e642334;
8'ha6 : rvCrc[30] <= 32'h6cf637bc;
8'ha7 : rvCrc[30] <= 32'h4d783bc4;
8'ha8 : rvCrc[30] <= 32'ha16360db;
8'ha9 : rvCrc[30] <= 32'h80ed6ca3;
8'haa : rvCrc[30] <= 32'he27f782b;
8'hab : rvCrc[30] <= 32'hc3f17453;
8'hac : rvCrc[30] <= 32'h275b513b;
8'had : rvCrc[30] <= 32'h06d55d43;
8'hae : rvCrc[30] <= 32'h644749cb;
8'haf : rvCrc[30] <= 32'h45c945b3;
8'hb0 : rvCrc[30] <= 32'hb8b0e242;
8'hb1 : rvCrc[30] <= 32'h993eee3a;
8'hb2 : rvCrc[30] <= 32'hfbacfab2;
8'hb3 : rvCrc[30] <= 32'hda22f6ca;
8'hb4 : rvCrc[30] <= 32'h3e88d3a2;
8'hb5 : rvCrc[30] <= 32'h1f06dfda;
8'hb6 : rvCrc[30] <= 32'h7d94cb52;
8'hb7 : rvCrc[30] <= 32'h5c1ac72a;
8'hb8 : rvCrc[30] <= 32'hb0019c35;
8'hb9 : rvCrc[30] <= 32'h918f904d;
8'hba : rvCrc[30] <= 32'hf31d84c5;
8'hbb : rvCrc[30] <= 32'hd29388bd;
8'hbc : rvCrc[30] <= 32'h3639add5;
8'hbd : rvCrc[30] <= 32'h17b7a1ad;
8'hbe : rvCrc[30] <= 32'h7525b525;
8'hbf : rvCrc[30] <= 32'h54abb95d;
8'hc0 : rvCrc[30] <= 32'hce9c14c8;
8'hc1 : rvCrc[30] <= 32'hef1218b0;
8'hc2 : rvCrc[30] <= 32'h8d800c38;
8'hc3 : rvCrc[30] <= 32'hac0e0040;
8'hc4 : rvCrc[30] <= 32'h48a42528;
8'hc5 : rvCrc[30] <= 32'h692a2950;
8'hc6 : rvCrc[30] <= 32'h0bb83dd8;
8'hc7 : rvCrc[30] <= 32'h2a3631a0;
8'hc8 : rvCrc[30] <= 32'hc62d6abf;
8'hc9 : rvCrc[30] <= 32'he7a366c7;
8'hca : rvCrc[30] <= 32'h8531724f;
8'hcb : rvCrc[30] <= 32'ha4bf7e37;
8'hcc : rvCrc[30] <= 32'h40155b5f;
8'hcd : rvCrc[30] <= 32'h619b5727;
8'hce : rvCrc[30] <= 32'h030943af;
8'hcf : rvCrc[30] <= 32'h22874fd7;
8'hd0 : rvCrc[30] <= 32'hdffee826;
8'hd1 : rvCrc[30] <= 32'hfe70e45e;
8'hd2 : rvCrc[30] <= 32'h9ce2f0d6;
8'hd3 : rvCrc[30] <= 32'hbd6cfcae;
8'hd4 : rvCrc[30] <= 32'h59c6d9c6;
8'hd5 : rvCrc[30] <= 32'h7848d5be;
8'hd6 : rvCrc[30] <= 32'h1adac136;
8'hd7 : rvCrc[30] <= 32'h3b54cd4e;
8'hd8 : rvCrc[30] <= 32'hd74f9651;
8'hd9 : rvCrc[30] <= 32'hf6c19a29;
8'hda : rvCrc[30] <= 32'h94538ea1;
8'hdb : rvCrc[30] <= 32'hb5dd82d9;
8'hdc : rvCrc[30] <= 32'h5177a7b1;
8'hdd : rvCrc[30] <= 32'h70f9abc9;
8'hde : rvCrc[30] <= 32'h126bbf41;
8'hdf : rvCrc[30] <= 32'h33e5b339;
8'he0 : rvCrc[30] <= 32'hec59ed14;
8'he1 : rvCrc[30] <= 32'hcdd7e16c;
8'he2 : rvCrc[30] <= 32'haf45f5e4;
8'he3 : rvCrc[30] <= 32'h8ecbf99c;
8'he4 : rvCrc[30] <= 32'h6a61dcf4;
8'he5 : rvCrc[30] <= 32'h4befd08c;
8'he6 : rvCrc[30] <= 32'h297dc404;
8'he7 : rvCrc[30] <= 32'h08f3c87c;
8'he8 : rvCrc[30] <= 32'he4e89363;
8'he9 : rvCrc[30] <= 32'hc5669f1b;
8'hea : rvCrc[30] <= 32'ha7f48b93;
8'heb : rvCrc[30] <= 32'h867a87eb;
8'hec : rvCrc[30] <= 32'h62d0a283;
8'hed : rvCrc[30] <= 32'h435eaefb;
8'hee : rvCrc[30] <= 32'h21ccba73;
8'hef : rvCrc[30] <= 32'h0042b60b;
8'hf0 : rvCrc[30] <= 32'hfd3b11fa;
8'hf1 : rvCrc[30] <= 32'hdcb51d82;
8'hf2 : rvCrc[30] <= 32'hbe27090a;
8'hf3 : rvCrc[30] <= 32'h9fa90572;
8'hf4 : rvCrc[30] <= 32'h7b03201a;
8'hf5 : rvCrc[30] <= 32'h5a8d2c62;
8'hf6 : rvCrc[30] <= 32'h381f38ea;
8'hf7 : rvCrc[30] <= 32'h19913492;
8'hf8 : rvCrc[30] <= 32'hf58a6f8d;
8'hf9 : rvCrc[30] <= 32'hd40463f5;
8'hfa : rvCrc[30] <= 32'hb696777d;
8'hfb : rvCrc[30] <= 32'h97187b05;
8'hfc : rvCrc[30] <= 32'h73b25e6d;
8'hfd : rvCrc[30] <= 32'h523c5215;
8'hfe : rvCrc[30] <= 32'h30ae469d;
8'hff : rvCrc[30] <= 32'h11204ae5;
endcase
case(iv_Input[255:248])
8'h00 : rvCrc[31] <= 32'h00000000;
8'h01 : rvCrc[31] <= 32'h12eed357;
8'h02 : rvCrc[31] <= 32'h25dda6ae;
8'h03 : rvCrc[31] <= 32'h373375f9;
8'h04 : rvCrc[31] <= 32'h4bbb4d5c;
8'h05 : rvCrc[31] <= 32'h59559e0b;
8'h06 : rvCrc[31] <= 32'h6e66ebf2;
8'h07 : rvCrc[31] <= 32'h7c8838a5;
8'h08 : rvCrc[31] <= 32'h97769ab8;
8'h09 : rvCrc[31] <= 32'h859849ef;
8'h0a : rvCrc[31] <= 32'hb2ab3c16;
8'h0b : rvCrc[31] <= 32'ha045ef41;
8'h0c : rvCrc[31] <= 32'hdccdd7e4;
8'h0d : rvCrc[31] <= 32'hce2304b3;
8'h0e : rvCrc[31] <= 32'hf910714a;
8'h0f : rvCrc[31] <= 32'hebfea21d;
8'h10 : rvCrc[31] <= 32'h2a2c28c7;
8'h11 : rvCrc[31] <= 32'h38c2fb90;
8'h12 : rvCrc[31] <= 32'h0ff18e69;
8'h13 : rvCrc[31] <= 32'h1d1f5d3e;
8'h14 : rvCrc[31] <= 32'h6197659b;
8'h15 : rvCrc[31] <= 32'h7379b6cc;
8'h16 : rvCrc[31] <= 32'h444ac335;
8'h17 : rvCrc[31] <= 32'h56a41062;
8'h18 : rvCrc[31] <= 32'hbd5ab27f;
8'h19 : rvCrc[31] <= 32'hafb46128;
8'h1a : rvCrc[31] <= 32'h988714d1;
8'h1b : rvCrc[31] <= 32'h8a69c786;
8'h1c : rvCrc[31] <= 32'hf6e1ff23;
8'h1d : rvCrc[31] <= 32'he40f2c74;
8'h1e : rvCrc[31] <= 32'hd33c598d;
8'h1f : rvCrc[31] <= 32'hc1d28ada;
8'h20 : rvCrc[31] <= 32'h5458518e;
8'h21 : rvCrc[31] <= 32'h46b682d9;
8'h22 : rvCrc[31] <= 32'h7185f720;
8'h23 : rvCrc[31] <= 32'h636b2477;
8'h24 : rvCrc[31] <= 32'h1fe31cd2;
8'h25 : rvCrc[31] <= 32'h0d0dcf85;
8'h26 : rvCrc[31] <= 32'h3a3eba7c;
8'h27 : rvCrc[31] <= 32'h28d0692b;
8'h28 : rvCrc[31] <= 32'hc32ecb36;
8'h29 : rvCrc[31] <= 32'hd1c01861;
8'h2a : rvCrc[31] <= 32'he6f36d98;
8'h2b : rvCrc[31] <= 32'hf41dbecf;
8'h2c : rvCrc[31] <= 32'h8895866a;
8'h2d : rvCrc[31] <= 32'h9a7b553d;
8'h2e : rvCrc[31] <= 32'had4820c4;
8'h2f : rvCrc[31] <= 32'hbfa6f393;
8'h30 : rvCrc[31] <= 32'h7e747949;
8'h31 : rvCrc[31] <= 32'h6c9aaa1e;
8'h32 : rvCrc[31] <= 32'h5ba9dfe7;
8'h33 : rvCrc[31] <= 32'h49470cb0;
8'h34 : rvCrc[31] <= 32'h35cf3415;
8'h35 : rvCrc[31] <= 32'h2721e742;
8'h36 : rvCrc[31] <= 32'h101292bb;
8'h37 : rvCrc[31] <= 32'h02fc41ec;
8'h38 : rvCrc[31] <= 32'he902e3f1;
8'h39 : rvCrc[31] <= 32'hfbec30a6;
8'h3a : rvCrc[31] <= 32'hccdf455f;
8'h3b : rvCrc[31] <= 32'hde319608;
8'h3c : rvCrc[31] <= 32'ha2b9aead;
8'h3d : rvCrc[31] <= 32'hb0577dfa;
8'h3e : rvCrc[31] <= 32'h87640803;
8'h3f : rvCrc[31] <= 32'h958adb54;
8'h40 : rvCrc[31] <= 32'ha8b0a31c;
8'h41 : rvCrc[31] <= 32'hba5e704b;
8'h42 : rvCrc[31] <= 32'h8d6d05b2;
8'h43 : rvCrc[31] <= 32'h9f83d6e5;
8'h44 : rvCrc[31] <= 32'he30bee40;
8'h45 : rvCrc[31] <= 32'hf1e53d17;
8'h46 : rvCrc[31] <= 32'hc6d648ee;
8'h47 : rvCrc[31] <= 32'hd4389bb9;
8'h48 : rvCrc[31] <= 32'h3fc639a4;
8'h49 : rvCrc[31] <= 32'h2d28eaf3;
8'h4a : rvCrc[31] <= 32'h1a1b9f0a;
8'h4b : rvCrc[31] <= 32'h08f54c5d;
8'h4c : rvCrc[31] <= 32'h747d74f8;
8'h4d : rvCrc[31] <= 32'h6693a7af;
8'h4e : rvCrc[31] <= 32'h51a0d256;
8'h4f : rvCrc[31] <= 32'h434e0101;
8'h50 : rvCrc[31] <= 32'h829c8bdb;
8'h51 : rvCrc[31] <= 32'h9072588c;
8'h52 : rvCrc[31] <= 32'ha7412d75;
8'h53 : rvCrc[31] <= 32'hb5affe22;
8'h54 : rvCrc[31] <= 32'hc927c687;
8'h55 : rvCrc[31] <= 32'hdbc915d0;
8'h56 : rvCrc[31] <= 32'hecfa6029;
8'h57 : rvCrc[31] <= 32'hfe14b37e;
8'h58 : rvCrc[31] <= 32'h15ea1163;
8'h59 : rvCrc[31] <= 32'h0704c234;
8'h5a : rvCrc[31] <= 32'h3037b7cd;
8'h5b : rvCrc[31] <= 32'h22d9649a;
8'h5c : rvCrc[31] <= 32'h5e515c3f;
8'h5d : rvCrc[31] <= 32'h4cbf8f68;
8'h5e : rvCrc[31] <= 32'h7b8cfa91;
8'h5f : rvCrc[31] <= 32'h696229c6;
8'h60 : rvCrc[31] <= 32'hfce8f292;
8'h61 : rvCrc[31] <= 32'hee0621c5;
8'h62 : rvCrc[31] <= 32'hd935543c;
8'h63 : rvCrc[31] <= 32'hcbdb876b;
8'h64 : rvCrc[31] <= 32'hb753bfce;
8'h65 : rvCrc[31] <= 32'ha5bd6c99;
8'h66 : rvCrc[31] <= 32'h928e1960;
8'h67 : rvCrc[31] <= 32'h8060ca37;
8'h68 : rvCrc[31] <= 32'h6b9e682a;
8'h69 : rvCrc[31] <= 32'h7970bb7d;
8'h6a : rvCrc[31] <= 32'h4e43ce84;
8'h6b : rvCrc[31] <= 32'h5cad1dd3;
8'h6c : rvCrc[31] <= 32'h20252576;
8'h6d : rvCrc[31] <= 32'h32cbf621;
8'h6e : rvCrc[31] <= 32'h05f883d8;
8'h6f : rvCrc[31] <= 32'h1716508f;
8'h70 : rvCrc[31] <= 32'hd6c4da55;
8'h71 : rvCrc[31] <= 32'hc42a0902;
8'h72 : rvCrc[31] <= 32'hf3197cfb;
8'h73 : rvCrc[31] <= 32'he1f7afac;
8'h74 : rvCrc[31] <= 32'h9d7f9709;
8'h75 : rvCrc[31] <= 32'h8f91445e;
8'h76 : rvCrc[31] <= 32'hb8a231a7;
8'h77 : rvCrc[31] <= 32'haa4ce2f0;
8'h78 : rvCrc[31] <= 32'h41b240ed;
8'h79 : rvCrc[31] <= 32'h535c93ba;
8'h7a : rvCrc[31] <= 32'h646fe643;
8'h7b : rvCrc[31] <= 32'h76813514;
8'h7c : rvCrc[31] <= 32'h0a090db1;
8'h7d : rvCrc[31] <= 32'h18e7dee6;
8'h7e : rvCrc[31] <= 32'h2fd4ab1f;
8'h7f : rvCrc[31] <= 32'h3d3a7848;
8'h80 : rvCrc[31] <= 32'h55a05b8f;
8'h81 : rvCrc[31] <= 32'h474e88d8;
8'h82 : rvCrc[31] <= 32'h707dfd21;
8'h83 : rvCrc[31] <= 32'h62932e76;
8'h84 : rvCrc[31] <= 32'h1e1b16d3;
8'h85 : rvCrc[31] <= 32'h0cf5c584;
8'h86 : rvCrc[31] <= 32'h3bc6b07d;
8'h87 : rvCrc[31] <= 32'h2928632a;
8'h88 : rvCrc[31] <= 32'hc2d6c137;
8'h89 : rvCrc[31] <= 32'hd0381260;
8'h8a : rvCrc[31] <= 32'he70b6799;
8'h8b : rvCrc[31] <= 32'hf5e5b4ce;
8'h8c : rvCrc[31] <= 32'h896d8c6b;
8'h8d : rvCrc[31] <= 32'h9b835f3c;
8'h8e : rvCrc[31] <= 32'hacb02ac5;
8'h8f : rvCrc[31] <= 32'hbe5ef992;
8'h90 : rvCrc[31] <= 32'h7f8c7348;
8'h91 : rvCrc[31] <= 32'h6d62a01f;
8'h92 : rvCrc[31] <= 32'h5a51d5e6;
8'h93 : rvCrc[31] <= 32'h48bf06b1;
8'h94 : rvCrc[31] <= 32'h34373e14;
8'h95 : rvCrc[31] <= 32'h26d9ed43;
8'h96 : rvCrc[31] <= 32'h11ea98ba;
8'h97 : rvCrc[31] <= 32'h03044bed;
8'h98 : rvCrc[31] <= 32'he8fae9f0;
8'h99 : rvCrc[31] <= 32'hfa143aa7;
8'h9a : rvCrc[31] <= 32'hcd274f5e;
8'h9b : rvCrc[31] <= 32'hdfc99c09;
8'h9c : rvCrc[31] <= 32'ha341a4ac;
8'h9d : rvCrc[31] <= 32'hb1af77fb;
8'h9e : rvCrc[31] <= 32'h869c0202;
8'h9f : rvCrc[31] <= 32'h9472d155;
8'ha0 : rvCrc[31] <= 32'h01f80a01;
8'ha1 : rvCrc[31] <= 32'h1316d956;
8'ha2 : rvCrc[31] <= 32'h2425acaf;
8'ha3 : rvCrc[31] <= 32'h36cb7ff8;
8'ha4 : rvCrc[31] <= 32'h4a43475d;
8'ha5 : rvCrc[31] <= 32'h58ad940a;
8'ha6 : rvCrc[31] <= 32'h6f9ee1f3;
8'ha7 : rvCrc[31] <= 32'h7d7032a4;
8'ha8 : rvCrc[31] <= 32'h968e90b9;
8'ha9 : rvCrc[31] <= 32'h846043ee;
8'haa : rvCrc[31] <= 32'hb3533617;
8'hab : rvCrc[31] <= 32'ha1bde540;
8'hac : rvCrc[31] <= 32'hdd35dde5;
8'had : rvCrc[31] <= 32'hcfdb0eb2;
8'hae : rvCrc[31] <= 32'hf8e87b4b;
8'haf : rvCrc[31] <= 32'hea06a81c;
8'hb0 : rvCrc[31] <= 32'h2bd422c6;
8'hb1 : rvCrc[31] <= 32'h393af191;
8'hb2 : rvCrc[31] <= 32'h0e098468;
8'hb3 : rvCrc[31] <= 32'h1ce7573f;
8'hb4 : rvCrc[31] <= 32'h606f6f9a;
8'hb5 : rvCrc[31] <= 32'h7281bccd;
8'hb6 : rvCrc[31] <= 32'h45b2c934;
8'hb7 : rvCrc[31] <= 32'h575c1a63;
8'hb8 : rvCrc[31] <= 32'hbca2b87e;
8'hb9 : rvCrc[31] <= 32'hae4c6b29;
8'hba : rvCrc[31] <= 32'h997f1ed0;
8'hbb : rvCrc[31] <= 32'h8b91cd87;
8'hbc : rvCrc[31] <= 32'hf719f522;
8'hbd : rvCrc[31] <= 32'he5f72675;
8'hbe : rvCrc[31] <= 32'hd2c4538c;
8'hbf : rvCrc[31] <= 32'hc02a80db;
8'hc0 : rvCrc[31] <= 32'hfd10f893;
8'hc1 : rvCrc[31] <= 32'heffe2bc4;
8'hc2 : rvCrc[31] <= 32'hd8cd5e3d;
8'hc3 : rvCrc[31] <= 32'hca238d6a;
8'hc4 : rvCrc[31] <= 32'hb6abb5cf;
8'hc5 : rvCrc[31] <= 32'ha4456698;
8'hc6 : rvCrc[31] <= 32'h93761361;
8'hc7 : rvCrc[31] <= 32'h8198c036;
8'hc8 : rvCrc[31] <= 32'h6a66622b;
8'hc9 : rvCrc[31] <= 32'h7888b17c;
8'hca : rvCrc[31] <= 32'h4fbbc485;
8'hcb : rvCrc[31] <= 32'h5d5517d2;
8'hcc : rvCrc[31] <= 32'h21dd2f77;
8'hcd : rvCrc[31] <= 32'h3333fc20;
8'hce : rvCrc[31] <= 32'h040089d9;
8'hcf : rvCrc[31] <= 32'h16ee5a8e;
8'hd0 : rvCrc[31] <= 32'hd73cd054;
8'hd1 : rvCrc[31] <= 32'hc5d20303;
8'hd2 : rvCrc[31] <= 32'hf2e176fa;
8'hd3 : rvCrc[31] <= 32'he00fa5ad;
8'hd4 : rvCrc[31] <= 32'h9c879d08;
8'hd5 : rvCrc[31] <= 32'h8e694e5f;
8'hd6 : rvCrc[31] <= 32'hb95a3ba6;
8'hd7 : rvCrc[31] <= 32'habb4e8f1;
8'hd8 : rvCrc[31] <= 32'h404a4aec;
8'hd9 : rvCrc[31] <= 32'h52a499bb;
8'hda : rvCrc[31] <= 32'h6597ec42;
8'hdb : rvCrc[31] <= 32'h77793f15;
8'hdc : rvCrc[31] <= 32'h0bf107b0;
8'hdd : rvCrc[31] <= 32'h191fd4e7;
8'hde : rvCrc[31] <= 32'h2e2ca11e;
8'hdf : rvCrc[31] <= 32'h3cc27249;
8'he0 : rvCrc[31] <= 32'ha948a91d;
8'he1 : rvCrc[31] <= 32'hbba67a4a;
8'he2 : rvCrc[31] <= 32'h8c950fb3;
8'he3 : rvCrc[31] <= 32'h9e7bdce4;
8'he4 : rvCrc[31] <= 32'he2f3e441;
8'he5 : rvCrc[31] <= 32'hf01d3716;
8'he6 : rvCrc[31] <= 32'hc72e42ef;
8'he7 : rvCrc[31] <= 32'hd5c091b8;
8'he8 : rvCrc[31] <= 32'h3e3e33a5;
8'he9 : rvCrc[31] <= 32'h2cd0e0f2;
8'hea : rvCrc[31] <= 32'h1be3950b;
8'heb : rvCrc[31] <= 32'h090d465c;
8'hec : rvCrc[31] <= 32'h75857ef9;
8'hed : rvCrc[31] <= 32'h676badae;
8'hee : rvCrc[31] <= 32'h5058d857;
8'hef : rvCrc[31] <= 32'h42b60b00;
8'hf0 : rvCrc[31] <= 32'h836481da;
8'hf1 : rvCrc[31] <= 32'h918a528d;
8'hf2 : rvCrc[31] <= 32'ha6b92774;
8'hf3 : rvCrc[31] <= 32'hb457f423;
8'hf4 : rvCrc[31] <= 32'hc8dfcc86;
8'hf5 : rvCrc[31] <= 32'hda311fd1;
8'hf6 : rvCrc[31] <= 32'hed026a28;
8'hf7 : rvCrc[31] <= 32'hffecb97f;
8'hf8 : rvCrc[31] <= 32'h14121b62;
8'hf9 : rvCrc[31] <= 32'h06fcc835;
8'hfa : rvCrc[31] <= 32'h31cfbdcc;
8'hfb : rvCrc[31] <= 32'h23216e9b;
8'hfc : rvCrc[31] <= 32'h5fa9563e;
8'hfd : rvCrc[31] <= 32'h4d478569;
8'hfe : rvCrc[31] <= 32'h7a74f090;
8'hff : rvCrc[31] <= 32'h689a23c7;
endcase
end
assign o32_Crc = rvCrc[0]^rvCrc[1]^rvCrc[2]^rvCrc[3]^rvCrc[4]^rvCrc[5]^rvCrc[6]^rvCrc[7]^rvCrc[8]^rvCrc[9]^rvCrc[10]^rvCrc[11]^rvCrc[12]^rvCrc[13]^rvCrc[14]^rvCrc[15]^rvCrc[16]^rvCrc[17]^rvCrc[18]^rvCrc[19]^rvCrc[20]^rvCrc[21]^rvCrc[22]^rvCrc[23]^rvCrc[24]^rvCrc[25]^rvCrc[26]^rvCrc[27]^rvCrc[28]^rvCrc[29]^rvCrc[30]^rvCrc[31];

endmodule 




